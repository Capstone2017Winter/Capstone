--megafunction wizard: %Altera SOPC Builder%
--GENERATION: STANDARD
--VERSION: WM1.0


--Legal Notice: (C)2013 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity altpll_inst_pll_slave_arbitrator is 
        port (
              -- inputs:
                 signal altpll_inst_pll_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_clock_0_out_read : IN STD_LOGIC;
                 signal niosII_system_clock_0_out_write : IN STD_LOGIC;
                 signal niosII_system_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal altpll_inst_pll_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal altpll_inst_pll_slave_read : OUT STD_LOGIC;
                 signal altpll_inst_pll_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal altpll_inst_pll_slave_reset : OUT STD_LOGIC;
                 signal altpll_inst_pll_slave_write : OUT STD_LOGIC;
                 signal altpll_inst_pll_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_altpll_inst_pll_slave_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_clock_0_out_granted_altpll_inst_pll_slave : OUT STD_LOGIC;
                 signal niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave : OUT STD_LOGIC;
                 signal niosII_system_clock_0_out_read_data_valid_altpll_inst_pll_slave : OUT STD_LOGIC;
                 signal niosII_system_clock_0_out_requests_altpll_inst_pll_slave : OUT STD_LOGIC
              );
end entity altpll_inst_pll_slave_arbitrator;


architecture europa of altpll_inst_pll_slave_arbitrator is
                signal altpll_inst_pll_slave_allgrants :  STD_LOGIC;
                signal altpll_inst_pll_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal altpll_inst_pll_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal altpll_inst_pll_slave_any_continuerequest :  STD_LOGIC;
                signal altpll_inst_pll_slave_arb_counter_enable :  STD_LOGIC;
                signal altpll_inst_pll_slave_arb_share_counter :  STD_LOGIC;
                signal altpll_inst_pll_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal altpll_inst_pll_slave_arb_share_set_values :  STD_LOGIC;
                signal altpll_inst_pll_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal altpll_inst_pll_slave_begins_xfer :  STD_LOGIC;
                signal altpll_inst_pll_slave_end_xfer :  STD_LOGIC;
                signal altpll_inst_pll_slave_firsttransfer :  STD_LOGIC;
                signal altpll_inst_pll_slave_grant_vector :  STD_LOGIC;
                signal altpll_inst_pll_slave_in_a_read_cycle :  STD_LOGIC;
                signal altpll_inst_pll_slave_in_a_write_cycle :  STD_LOGIC;
                signal altpll_inst_pll_slave_master_qreq_vector :  STD_LOGIC;
                signal altpll_inst_pll_slave_non_bursting_master_requests :  STD_LOGIC;
                signal altpll_inst_pll_slave_reg_firsttransfer :  STD_LOGIC;
                signal altpll_inst_pll_slave_slavearbiterlockenable :  STD_LOGIC;
                signal altpll_inst_pll_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal altpll_inst_pll_slave_unreg_firsttransfer :  STD_LOGIC;
                signal altpll_inst_pll_slave_waits_for_read :  STD_LOGIC;
                signal altpll_inst_pll_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_altpll_inst_pll_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_clock_0_out_granted_altpll_inst_pll_slave :  STD_LOGIC;
                signal internal_niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave :  STD_LOGIC;
                signal internal_niosII_system_clock_0_out_requests_altpll_inst_pll_slave :  STD_LOGIC;
                signal niosII_system_clock_0_out_arbiterlock :  STD_LOGIC;
                signal niosII_system_clock_0_out_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_clock_0_out_continuerequest :  STD_LOGIC;
                signal niosII_system_clock_0_out_saved_grant_altpll_inst_pll_slave :  STD_LOGIC;
                signal shifted_address_to_altpll_inst_pll_slave_from_niosII_system_clock_0_out :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal wait_for_altpll_inst_pll_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT altpll_inst_pll_slave_end_xfer;
    end if;

  end process;

  altpll_inst_pll_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave);
  --assign altpll_inst_pll_slave_readdata_from_sa = altpll_inst_pll_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  altpll_inst_pll_slave_readdata_from_sa <= altpll_inst_pll_slave_readdata;
  internal_niosII_system_clock_0_out_requests_altpll_inst_pll_slave <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_clock_0_out_read OR niosII_system_clock_0_out_write)))))));
  --altpll_inst_pll_slave_arb_share_counter set values, which is an e_mux
  altpll_inst_pll_slave_arb_share_set_values <= std_logic'('1');
  --altpll_inst_pll_slave_non_bursting_master_requests mux, which is an e_mux
  altpll_inst_pll_slave_non_bursting_master_requests <= internal_niosII_system_clock_0_out_requests_altpll_inst_pll_slave;
  --altpll_inst_pll_slave_any_bursting_master_saved_grant mux, which is an e_mux
  altpll_inst_pll_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --altpll_inst_pll_slave_arb_share_counter_next_value assignment, which is an e_assign
  altpll_inst_pll_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(altpll_inst_pll_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_inst_pll_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(altpll_inst_pll_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_inst_pll_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --altpll_inst_pll_slave_allgrants all slave grants, which is an e_mux
  altpll_inst_pll_slave_allgrants <= altpll_inst_pll_slave_grant_vector;
  --altpll_inst_pll_slave_end_xfer assignment, which is an e_assign
  altpll_inst_pll_slave_end_xfer <= NOT ((altpll_inst_pll_slave_waits_for_read OR altpll_inst_pll_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_altpll_inst_pll_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_altpll_inst_pll_slave <= altpll_inst_pll_slave_end_xfer AND (((NOT altpll_inst_pll_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --altpll_inst_pll_slave_arb_share_counter arbitration counter enable, which is an e_assign
  altpll_inst_pll_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_altpll_inst_pll_slave AND altpll_inst_pll_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_altpll_inst_pll_slave AND NOT altpll_inst_pll_slave_non_bursting_master_requests));
  --altpll_inst_pll_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      altpll_inst_pll_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(altpll_inst_pll_slave_arb_counter_enable) = '1' then 
        altpll_inst_pll_slave_arb_share_counter <= altpll_inst_pll_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --altpll_inst_pll_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      altpll_inst_pll_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((altpll_inst_pll_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_altpll_inst_pll_slave)) OR ((end_xfer_arb_share_counter_term_altpll_inst_pll_slave AND NOT altpll_inst_pll_slave_non_bursting_master_requests)))) = '1' then 
        altpll_inst_pll_slave_slavearbiterlockenable <= altpll_inst_pll_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_clock_0/out altpll_inst/pll_slave arbiterlock, which is an e_assign
  niosII_system_clock_0_out_arbiterlock <= altpll_inst_pll_slave_slavearbiterlockenable AND niosII_system_clock_0_out_continuerequest;
  --altpll_inst_pll_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  altpll_inst_pll_slave_slavearbiterlockenable2 <= altpll_inst_pll_slave_arb_share_counter_next_value;
  --niosII_system_clock_0/out altpll_inst/pll_slave arbiterlock2, which is an e_assign
  niosII_system_clock_0_out_arbiterlock2 <= altpll_inst_pll_slave_slavearbiterlockenable2 AND niosII_system_clock_0_out_continuerequest;
  --altpll_inst_pll_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  altpll_inst_pll_slave_any_continuerequest <= std_logic'('1');
  --niosII_system_clock_0_out_continuerequest continued request, which is an e_assign
  niosII_system_clock_0_out_continuerequest <= std_logic'('1');
  internal_niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave <= internal_niosII_system_clock_0_out_requests_altpll_inst_pll_slave;
  --altpll_inst_pll_slave_writedata mux, which is an e_mux
  altpll_inst_pll_slave_writedata <= niosII_system_clock_0_out_writedata;
  --master is always granted when requested
  internal_niosII_system_clock_0_out_granted_altpll_inst_pll_slave <= internal_niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave;
  --niosII_system_clock_0/out saved-grant altpll_inst/pll_slave, which is an e_assign
  niosII_system_clock_0_out_saved_grant_altpll_inst_pll_slave <= internal_niosII_system_clock_0_out_requests_altpll_inst_pll_slave;
  --allow new arb cycle for altpll_inst/pll_slave, which is an e_assign
  altpll_inst_pll_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  altpll_inst_pll_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  altpll_inst_pll_slave_master_qreq_vector <= std_logic'('1');
  --~altpll_inst_pll_slave_reset assignment, which is an e_assign
  altpll_inst_pll_slave_reset <= NOT reset_n;
  --altpll_inst_pll_slave_firsttransfer first transaction, which is an e_assign
  altpll_inst_pll_slave_firsttransfer <= A_WE_StdLogic((std_logic'(altpll_inst_pll_slave_begins_xfer) = '1'), altpll_inst_pll_slave_unreg_firsttransfer, altpll_inst_pll_slave_reg_firsttransfer);
  --altpll_inst_pll_slave_unreg_firsttransfer first transaction, which is an e_assign
  altpll_inst_pll_slave_unreg_firsttransfer <= NOT ((altpll_inst_pll_slave_slavearbiterlockenable AND altpll_inst_pll_slave_any_continuerequest));
  --altpll_inst_pll_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      altpll_inst_pll_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(altpll_inst_pll_slave_begins_xfer) = '1' then 
        altpll_inst_pll_slave_reg_firsttransfer <= altpll_inst_pll_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --altpll_inst_pll_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  altpll_inst_pll_slave_beginbursttransfer_internal <= altpll_inst_pll_slave_begins_xfer;
  --altpll_inst_pll_slave_read assignment, which is an e_mux
  altpll_inst_pll_slave_read <= internal_niosII_system_clock_0_out_granted_altpll_inst_pll_slave AND niosII_system_clock_0_out_read;
  --altpll_inst_pll_slave_write assignment, which is an e_mux
  altpll_inst_pll_slave_write <= internal_niosII_system_clock_0_out_granted_altpll_inst_pll_slave AND niosII_system_clock_0_out_write;
  shifted_address_to_altpll_inst_pll_slave_from_niosII_system_clock_0_out <= niosII_system_clock_0_out_address_to_slave;
  --altpll_inst_pll_slave_address mux, which is an e_mux
  altpll_inst_pll_slave_address <= A_EXT (A_SRL(shifted_address_to_altpll_inst_pll_slave_from_niosII_system_clock_0_out,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_altpll_inst_pll_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_altpll_inst_pll_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_altpll_inst_pll_slave_end_xfer <= altpll_inst_pll_slave_end_xfer;
    end if;

  end process;

  --altpll_inst_pll_slave_waits_for_read in a cycle, which is an e_mux
  altpll_inst_pll_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_inst_pll_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --altpll_inst_pll_slave_in_a_read_cycle assignment, which is an e_assign
  altpll_inst_pll_slave_in_a_read_cycle <= internal_niosII_system_clock_0_out_granted_altpll_inst_pll_slave AND niosII_system_clock_0_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= altpll_inst_pll_slave_in_a_read_cycle;
  --altpll_inst_pll_slave_waits_for_write in a cycle, which is an e_mux
  altpll_inst_pll_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_inst_pll_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --altpll_inst_pll_slave_in_a_write_cycle assignment, which is an e_assign
  altpll_inst_pll_slave_in_a_write_cycle <= internal_niosII_system_clock_0_out_granted_altpll_inst_pll_slave AND niosII_system_clock_0_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= altpll_inst_pll_slave_in_a_write_cycle;
  wait_for_altpll_inst_pll_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  niosII_system_clock_0_out_granted_altpll_inst_pll_slave <= internal_niosII_system_clock_0_out_granted_altpll_inst_pll_slave;
  --vhdl renameroo for output signals
  niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave <= internal_niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave;
  --vhdl renameroo for output signals
  niosII_system_clock_0_out_requests_altpll_inst_pll_slave <= internal_niosII_system_clock_0_out_requests_altpll_inst_pll_slave;
--synthesis translate_off
    --altpll_inst/pll_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_jtag_debug_module_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_address_to_slave : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal niosII_system_burst_0_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_0_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_0_downstream_debugaccess : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_1_downstream_address_to_slave : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal niosII_system_burst_1_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_1_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_1_downstream_debugaccess : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal cpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_jtag_debug_module_reset_n : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_write : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_jtag_debug_module_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module : OUT STD_LOGIC
              );
end entity cpu_jtag_debug_module_arbitrator;


architecture europa of cpu_jtag_debug_module_arbitrator is
                signal cpu_jtag_debug_module_allgrants :  STD_LOGIC;
                signal cpu_jtag_debug_module_allow_new_arb_cycle :  STD_LOGIC;
                signal cpu_jtag_debug_module_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cpu_jtag_debug_module_any_continuerequest :  STD_LOGIC;
                signal cpu_jtag_debug_module_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_arb_counter_enable :  STD_LOGIC;
                signal cpu_jtag_debug_module_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_jtag_debug_module_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_jtag_debug_module_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_jtag_debug_module_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_arbitration_holdoff_internal :  STD_LOGIC;
                signal cpu_jtag_debug_module_beginbursttransfer_internal :  STD_LOGIC;
                signal cpu_jtag_debug_module_begins_xfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_jtag_debug_module_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_firsttransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_in_a_read_cycle :  STD_LOGIC;
                signal cpu_jtag_debug_module_in_a_write_cycle :  STD_LOGIC;
                signal cpu_jtag_debug_module_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_non_bursting_master_requests :  STD_LOGIC;
                signal cpu_jtag_debug_module_reg_firsttransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_slavearbiterlockenable :  STD_LOGIC;
                signal cpu_jtag_debug_module_slavearbiterlockenable2 :  STD_LOGIC;
                signal cpu_jtag_debug_module_unreg_firsttransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_waits_for_read :  STD_LOGIC;
                signal cpu_jtag_debug_module_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cpu_jtag_debug_module :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_niosII_system_burst_0_downstream_granted_slave_cpu_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_niosII_system_burst_1_downstream_granted_slave_cpu_jtag_debug_module :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_saved_grant_cpu_jtag_debug_module :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_saved_grant_cpu_jtag_debug_module :  STD_LOGIC;
                signal shifted_address_to_cpu_jtag_debug_module_from_niosII_system_burst_0_downstream :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal shifted_address_to_cpu_jtag_debug_module_from_niosII_system_burst_1_downstream :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal wait_for_cpu_jtag_debug_module_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  cpu_jtag_debug_module_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module OR internal_niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module));
  --assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_jtag_debug_module_readdata_from_sa <= cpu_jtag_debug_module_readdata;
  internal_niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_0_downstream_read OR niosII_system_burst_0_downstream_write)))))));
  --cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  cpu_jtag_debug_module_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_0_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_1_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_0_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_1_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001"))))), 4);
  --cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  cpu_jtag_debug_module_non_bursting_master_requests <= std_logic'('0');
  --cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  cpu_jtag_debug_module_any_bursting_master_saved_grant <= ((niosII_system_burst_0_downstream_saved_grant_cpu_jtag_debug_module OR niosII_system_burst_1_downstream_saved_grant_cpu_jtag_debug_module) OR niosII_system_burst_0_downstream_saved_grant_cpu_jtag_debug_module) OR niosII_system_burst_1_downstream_saved_grant_cpu_jtag_debug_module;
  --cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  cpu_jtag_debug_module_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(cpu_jtag_debug_module_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (cpu_jtag_debug_module_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(cpu_jtag_debug_module_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (cpu_jtag_debug_module_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  cpu_jtag_debug_module_allgrants <= (((or_reduce(cpu_jtag_debug_module_grant_vector)) OR (or_reduce(cpu_jtag_debug_module_grant_vector))) OR (or_reduce(cpu_jtag_debug_module_grant_vector))) OR (or_reduce(cpu_jtag_debug_module_grant_vector));
  --cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  cpu_jtag_debug_module_end_xfer <= NOT ((cpu_jtag_debug_module_waits_for_read OR cpu_jtag_debug_module_waits_for_write));
  --end_xfer_arb_share_counter_term_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cpu_jtag_debug_module <= cpu_jtag_debug_module_end_xfer AND (((NOT cpu_jtag_debug_module_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  cpu_jtag_debug_module_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cpu_jtag_debug_module AND cpu_jtag_debug_module_allgrants)) OR ((end_xfer_arb_share_counter_term_cpu_jtag_debug_module AND NOT cpu_jtag_debug_module_non_bursting_master_requests));
  --cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_jtag_debug_module_arb_counter_enable) = '1' then 
        cpu_jtag_debug_module_arb_share_counter <= cpu_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(cpu_jtag_debug_module_master_qreq_vector) AND end_xfer_arb_share_counter_term_cpu_jtag_debug_module)) OR ((end_xfer_arb_share_counter_term_cpu_jtag_debug_module AND NOT cpu_jtag_debug_module_non_bursting_master_requests)))) = '1' then 
        cpu_jtag_debug_module_slavearbiterlockenable <= or_reduce(cpu_jtag_debug_module_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_0/downstream cpu/jtag_debug_module arbiterlock, which is an e_assign
  niosII_system_burst_0_downstream_arbiterlock <= cpu_jtag_debug_module_slavearbiterlockenable AND niosII_system_burst_0_downstream_continuerequest;
  --cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cpu_jtag_debug_module_slavearbiterlockenable2 <= or_reduce(cpu_jtag_debug_module_arb_share_counter_next_value);
  --niosII_system_burst_0/downstream cpu/jtag_debug_module arbiterlock2, which is an e_assign
  niosII_system_burst_0_downstream_arbiterlock2 <= cpu_jtag_debug_module_slavearbiterlockenable2 AND niosII_system_burst_0_downstream_continuerequest;
  --niosII_system_burst_1/downstream cpu/jtag_debug_module arbiterlock, which is an e_assign
  niosII_system_burst_1_downstream_arbiterlock <= cpu_jtag_debug_module_slavearbiterlockenable AND niosII_system_burst_1_downstream_continuerequest;
  --niosII_system_burst_1/downstream cpu/jtag_debug_module arbiterlock2, which is an e_assign
  niosII_system_burst_1_downstream_arbiterlock2 <= cpu_jtag_debug_module_slavearbiterlockenable2 AND niosII_system_burst_1_downstream_continuerequest;
  --niosII_system_burst_1/downstream granted cpu/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_niosII_system_burst_1_downstream_granted_slave_cpu_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_niosII_system_burst_1_downstream_granted_slave_cpu_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(niosII_system_burst_1_downstream_saved_grant_cpu_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_1_downstream_granted_slave_cpu_jtag_debug_module))))));
    end if;

  end process;

  --niosII_system_burst_1_downstream_continuerequest continued request, which is an e_mux
  niosII_system_burst_1_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_1_downstream_granted_slave_cpu_jtag_debug_module))) AND std_logic_vector'("00000000000000000000000000000001")));
  --cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  cpu_jtag_debug_module_any_continuerequest <= niosII_system_burst_1_downstream_continuerequest OR niosII_system_burst_0_downstream_continuerequest;
  internal_niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module <= internal_niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module AND NOT ((((niosII_system_burst_0_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_0_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR niosII_system_burst_1_downstream_arbiterlock));
  --local readdatavalid niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module <= (internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module AND niosII_system_burst_0_downstream_read) AND NOT cpu_jtag_debug_module_waits_for_read;
  --cpu_jtag_debug_module_writedata mux, which is an e_mux
  cpu_jtag_debug_module_writedata <= A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module)) = '1'), niosII_system_burst_0_downstream_writedata, niosII_system_burst_1_downstream_writedata);
  internal_niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_1_downstream_read OR niosII_system_burst_1_downstream_write)))))));
  --niosII_system_burst_0/downstream granted cpu/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_niosII_system_burst_0_downstream_granted_slave_cpu_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_niosII_system_burst_0_downstream_granted_slave_cpu_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(niosII_system_burst_0_downstream_saved_grant_cpu_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_0_downstream_granted_slave_cpu_jtag_debug_module))))));
    end if;

  end process;

  --niosII_system_burst_0_downstream_continuerequest continued request, which is an e_mux
  niosII_system_burst_0_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_0_downstream_granted_slave_cpu_jtag_debug_module))) AND std_logic_vector'("00000000000000000000000000000001")));
  internal_niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module <= internal_niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module AND NOT ((((niosII_system_burst_1_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_1_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR niosII_system_burst_0_downstream_arbiterlock));
  --local readdatavalid niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module <= (internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module AND niosII_system_burst_1_downstream_read) AND NOT cpu_jtag_debug_module_waits_for_read;
  --allow new arb cycle for cpu/jtag_debug_module, which is an e_assign
  cpu_jtag_debug_module_allow_new_arb_cycle <= NOT niosII_system_burst_0_downstream_arbiterlock AND NOT niosII_system_burst_1_downstream_arbiterlock;
  --niosII_system_burst_1/downstream assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  cpu_jtag_debug_module_master_qreq_vector(0) <= internal_niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module;
  --niosII_system_burst_1/downstream grant cpu/jtag_debug_module, which is an e_assign
  internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module <= cpu_jtag_debug_module_grant_vector(0);
  --niosII_system_burst_1/downstream saved-grant cpu/jtag_debug_module, which is an e_assign
  niosII_system_burst_1_downstream_saved_grant_cpu_jtag_debug_module <= cpu_jtag_debug_module_arb_winner(0);
  --niosII_system_burst_0/downstream assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  cpu_jtag_debug_module_master_qreq_vector(1) <= internal_niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module;
  --niosII_system_burst_0/downstream grant cpu/jtag_debug_module, which is an e_assign
  internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module <= cpu_jtag_debug_module_grant_vector(1);
  --niosII_system_burst_0/downstream saved-grant cpu/jtag_debug_module, which is an e_assign
  niosII_system_burst_0_downstream_saved_grant_cpu_jtag_debug_module <= cpu_jtag_debug_module_arb_winner(1);
  --cpu/jtag_debug_module chosen-master double-vector, which is an e_assign
  cpu_jtag_debug_module_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((cpu_jtag_debug_module_master_qreq_vector & cpu_jtag_debug_module_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT cpu_jtag_debug_module_master_qreq_vector & NOT cpu_jtag_debug_module_master_qreq_vector))) + (std_logic_vector'("000") & (cpu_jtag_debug_module_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  cpu_jtag_debug_module_arb_winner <= A_WE_StdLogicVector((std_logic'(((cpu_jtag_debug_module_allow_new_arb_cycle AND or_reduce(cpu_jtag_debug_module_grant_vector)))) = '1'), cpu_jtag_debug_module_grant_vector, cpu_jtag_debug_module_saved_chosen_master_vector);
  --saved cpu_jtag_debug_module_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_jtag_debug_module_allow_new_arb_cycle) = '1' then 
        cpu_jtag_debug_module_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(cpu_jtag_debug_module_grant_vector)) = '1'), cpu_jtag_debug_module_grant_vector, cpu_jtag_debug_module_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  cpu_jtag_debug_module_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((cpu_jtag_debug_module_chosen_master_double_vector(1) OR cpu_jtag_debug_module_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((cpu_jtag_debug_module_chosen_master_double_vector(0) OR cpu_jtag_debug_module_chosen_master_double_vector(2)))));
  --cpu/jtag_debug_module chosen master rotated left, which is an e_assign
  cpu_jtag_debug_module_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(cpu_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(cpu_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --cpu/jtag_debug_module's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(cpu_jtag_debug_module_grant_vector)) = '1' then 
        cpu_jtag_debug_module_arb_addend <= A_WE_StdLogicVector((std_logic'(cpu_jtag_debug_module_end_xfer) = '1'), cpu_jtag_debug_module_chosen_master_rot_left, cpu_jtag_debug_module_grant_vector);
      end if;
    end if;

  end process;

  cpu_jtag_debug_module_begintransfer <= cpu_jtag_debug_module_begins_xfer;
  --cpu_jtag_debug_module_reset_n assignment, which is an e_assign
  cpu_jtag_debug_module_reset_n <= reset_n;
  --assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_jtag_debug_module_resetrequest_from_sa <= cpu_jtag_debug_module_resetrequest;
  cpu_jtag_debug_module_chipselect <= internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module OR internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module;
  --cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  cpu_jtag_debug_module_firsttransfer <= A_WE_StdLogic((std_logic'(cpu_jtag_debug_module_begins_xfer) = '1'), cpu_jtag_debug_module_unreg_firsttransfer, cpu_jtag_debug_module_reg_firsttransfer);
  --cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  cpu_jtag_debug_module_unreg_firsttransfer <= NOT ((cpu_jtag_debug_module_slavearbiterlockenable AND cpu_jtag_debug_module_any_continuerequest));
  --cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_jtag_debug_module_begins_xfer) = '1' then 
        cpu_jtag_debug_module_reg_firsttransfer <= cpu_jtag_debug_module_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cpu_jtag_debug_module_beginbursttransfer_internal <= cpu_jtag_debug_module_begins_xfer;
  --cpu_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  cpu_jtag_debug_module_arbitration_holdoff_internal <= cpu_jtag_debug_module_begins_xfer AND cpu_jtag_debug_module_firsttransfer;
  --cpu_jtag_debug_module_write assignment, which is an e_mux
  cpu_jtag_debug_module_write <= ((internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module AND niosII_system_burst_0_downstream_write)) OR ((internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module AND niosII_system_burst_1_downstream_write));
  shifted_address_to_cpu_jtag_debug_module_from_niosII_system_burst_0_downstream <= niosII_system_burst_0_downstream_address_to_slave;
  --cpu_jtag_debug_module_address mux, which is an e_mux
  cpu_jtag_debug_module_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module)) = '1'), (A_SRL(shifted_address_to_cpu_jtag_debug_module_from_niosII_system_burst_0_downstream,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_cpu_jtag_debug_module_from_niosII_system_burst_1_downstream,std_logic_vector'("00000000000000000000000000000010")))), 9);
  shifted_address_to_cpu_jtag_debug_module_from_niosII_system_burst_1_downstream <= niosII_system_burst_1_downstream_address_to_slave;
  --d1_cpu_jtag_debug_module_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cpu_jtag_debug_module_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cpu_jtag_debug_module_end_xfer <= cpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  --cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  cpu_jtag_debug_module_waits_for_read <= cpu_jtag_debug_module_in_a_read_cycle AND cpu_jtag_debug_module_begins_xfer;
  --cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  cpu_jtag_debug_module_in_a_read_cycle <= ((internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module AND niosII_system_burst_0_downstream_read)) OR ((internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module AND niosII_system_burst_1_downstream_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cpu_jtag_debug_module_in_a_read_cycle;
  --cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  cpu_jtag_debug_module_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  cpu_jtag_debug_module_in_a_write_cycle <= ((internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module AND niosII_system_burst_0_downstream_write)) OR ((internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module AND niosII_system_burst_1_downstream_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cpu_jtag_debug_module_in_a_write_cycle;
  wait_for_cpu_jtag_debug_module_counter <= std_logic'('0');
  --cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  cpu_jtag_debug_module_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_0_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_1_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  --debugaccess mux, which is an e_mux
  cpu_jtag_debug_module_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_0_downstream_debugaccess))), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_1_downstream_debugaccess))), std_logic_vector'("00000000000000000000000000000000"))));
  --vhdl renameroo for output signals
  niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module <= internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module <= internal_niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module <= internal_niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module <= internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module <= internal_niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module <= internal_niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module;
--synthesis translate_off
    --cpu/jtag_debug_module enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_0/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_0_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line, now);
          write(write_line, string'(": "));
          write(write_line, string'("niosII_system_burst_0/downstream drove 0 on its 'arbitrationshare' port while accessing slave cpu/jtag_debug_module"));
          write(output, write_line.all);
          deallocate (write_line);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_0/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line1 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_0_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line1, now);
          write(write_line1, string'(": "));
          write(write_line1, string'("niosII_system_burst_0/downstream drove 0 on its 'burstcount' port while accessing slave cpu/jtag_debug_module"));
          write(output, write_line1.all);
          deallocate (write_line1);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_1/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line2 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_1_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line2, now);
          write(write_line2, string'(": "));
          write(write_line2, string'("niosII_system_burst_1/downstream drove 0 on its 'arbitrationshare' port while accessing slave cpu/jtag_debug_module"));
          write(output, write_line2.all);
          deallocate (write_line2);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_1/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line3 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_1_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line3, now);
          write(write_line3, string'(": "));
          write(write_line3, string'("niosII_system_burst_1/downstream drove 0 on its 'burstcount' port while accessing slave cpu/jtag_debug_module"));
          write(output, write_line3.all);
          deallocate (write_line3);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line4 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line4, now);
          write(write_line4, string'(": "));
          write(write_line4, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line4.all);
          deallocate (write_line4);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line5 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(niosII_system_burst_0_downstream_saved_grant_cpu_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(niosII_system_burst_1_downstream_saved_grant_cpu_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line5, now);
          write(write_line5, string'(": "));
          write(write_line5, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line5.all);
          deallocate (write_line5);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_data_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable_niosII_system_burst_11_upstream : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_byteenable_niosII_system_burst_13_upstream : IN STD_LOGIC;
                 signal cpu_data_master_byteenable_niosII_system_burst_20_upstream : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_granted_niosII_system_burst_11_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_13_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_14_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_15_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_16_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_17_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_18_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_1_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_20_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_21_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_3_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_4_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_5_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_6_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_7_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_8_upstream : IN STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_9_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_11_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_13_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_14_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_15_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_16_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_17_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_18_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_1_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_20_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_21_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_3_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_4_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_5_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_6_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_7_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_8_upstream : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_9_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_11_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_13_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_14_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_15_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_16_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_17_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_18_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_1_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_20_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_21_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_3_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_4_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_5_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_6_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_7_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_8_upstream : IN STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_9_upstream : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_niosII_system_burst_11_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_13_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_14_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_15_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_16_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_17_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_18_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_1_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_20_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_21_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_3_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_4_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_5_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_6_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_7_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_8_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_9_upstream_end_xfer : IN STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_irq_from_sa : IN STD_LOGIC;
                 signal high_res_timer_s1_irq_from_sa : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_11_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_11_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_13_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_13_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_14_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_14_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_15_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_15_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_16_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_16_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_17_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_17_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_18_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_18_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_1_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_1_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_20_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_20_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_21_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_21_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_3_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_3_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_4_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_4_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_5_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_5_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_6_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_6_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_7_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_7_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_8_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_8_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_9_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_9_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_timer_s1_irq_from_sa : IN STD_LOGIC;
                 signal uart_0_s1_irq_from_sa : IN STD_LOGIC;
                 signal uart_1_s1_irq_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal cpu_data_master_dbs_write_8 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal cpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_data_master_latency_counter : OUT STD_LOGIC;
                 signal cpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_data_master_readdatavalid : OUT STD_LOGIC;
                 signal cpu_data_master_waitrequest : OUT STD_LOGIC
              );
end entity cpu_data_master_arbitrator;


architecture europa of cpu_data_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpu_data_master_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_data_master_burstcount_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_data_master_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_data_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_is_granted_some_slave :  STD_LOGIC;
                signal cpu_data_master_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_read_but_no_slave_selected :  STD_LOGIC;
                signal cpu_data_master_read_last_time :  STD_LOGIC;
                signal cpu_data_master_run :  STD_LOGIC;
                signal cpu_data_master_write_last_time :  STD_LOGIC;
                signal cpu_data_master_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_latent_8_reg_segment_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_latent_8_reg_segment_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_latent_8_reg_segment_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_cpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_cpu_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_data_master_latency_counter :  STD_LOGIC;
                signal internal_cpu_data_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_cpu_data_master_latency_counter :  STD_LOGIC;
                signal p1_dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_dbs_latent_8_reg_segment_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_dbs_latent_8_reg_segment_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_dbs_latent_8_reg_segment_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_cpu_data_master_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_1_upstream OR NOT cpu_data_master_requests_niosII_system_burst_1_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_1_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_1_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_1_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_1_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_11_upstream OR NOT cpu_data_master_requests_niosII_system_burst_11_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_11_upstream OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_11_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_11_upstream OR NOT cpu_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_11_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_13_upstream OR NOT cpu_data_master_requests_niosII_system_burst_13_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_13_upstream OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_13_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_13_upstream OR NOT cpu_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_13_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((internal_cpu_data_master_dbs_address(1) AND internal_cpu_data_master_dbs_address(0))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_14_upstream OR NOT cpu_data_master_requests_niosII_system_burst_14_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_14_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_14_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_14_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_14_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_15_upstream OR NOT cpu_data_master_requests_niosII_system_burst_15_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_15_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_15_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_15_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_15_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_data_master_run <= ((r_0 AND r_1) AND r_2) AND r_3;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_16_upstream OR NOT cpu_data_master_requests_niosII_system_burst_16_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_16_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_16_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_16_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_16_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_17_upstream OR NOT cpu_data_master_requests_niosII_system_burst_17_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_17_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_17_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_17_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_17_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_18_upstream OR NOT cpu_data_master_requests_niosII_system_burst_18_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_18_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_18_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_18_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_18_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_20_upstream OR NOT cpu_data_master_requests_niosII_system_burst_20_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_20_upstream OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_20_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_20_upstream OR NOT cpu_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_20_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_21_upstream OR NOT cpu_data_master_requests_niosII_system_burst_21_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_21_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_21_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_21_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_21_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_3_upstream OR NOT cpu_data_master_requests_niosII_system_burst_3_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_3_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_3_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_3_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_3_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_4_upstream OR NOT cpu_data_master_requests_niosII_system_burst_4_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_4_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_4_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_4_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_4_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_5_upstream OR NOT cpu_data_master_requests_niosII_system_burst_5_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_5_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_5_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_5_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_5_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_6_upstream OR NOT cpu_data_master_requests_niosII_system_burst_6_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_6_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_6_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_6_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_6_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_7_upstream OR NOT cpu_data_master_requests_niosII_system_burst_7_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_7_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_7_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_7_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_7_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))));
  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_8_upstream OR NOT cpu_data_master_requests_niosII_system_burst_8_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_8_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_8_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_8_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_8_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_niosII_system_burst_9_upstream OR NOT cpu_data_master_requests_niosII_system_burst_9_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_9_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_9_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_niosII_system_burst_9_upstream OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_9_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))));
  --irq assign, which is an e_assign
  cpu_data_master_irq <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(uart_1_s1_irq_from_sa) & A_ToStdLogicVector(uart_0_s1_irq_from_sa) & A_ToStdLogicVector(dm9000a_inst_avalon_slave_0_irq_from_sa) & A_ToStdLogicVector(high_res_timer_s1_irq_from_sa) & A_ToStdLogicVector(sys_clk_timer_s1_irq_from_sa) & A_ToStdLogicVector(jtag_uart_avalon_jtag_slave_irq_from_sa));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_data_master_address_to_slave <= cpu_data_master_address(24 DOWNTO 0);
  --cpu_data_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_data_master_read_but_no_slave_selected <= (cpu_data_master_read AND cpu_data_master_run) AND NOT cpu_data_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  cpu_data_master_is_granted_some_slave <= (((((((((((((((cpu_data_master_granted_niosII_system_burst_1_upstream OR cpu_data_master_granted_niosII_system_burst_11_upstream) OR cpu_data_master_granted_niosII_system_burst_13_upstream) OR cpu_data_master_granted_niosII_system_burst_14_upstream) OR cpu_data_master_granted_niosII_system_burst_15_upstream) OR cpu_data_master_granted_niosII_system_burst_16_upstream) OR cpu_data_master_granted_niosII_system_burst_17_upstream) OR cpu_data_master_granted_niosII_system_burst_18_upstream) OR cpu_data_master_granted_niosII_system_burst_20_upstream) OR cpu_data_master_granted_niosII_system_burst_21_upstream) OR cpu_data_master_granted_niosII_system_burst_3_upstream) OR cpu_data_master_granted_niosII_system_burst_4_upstream) OR cpu_data_master_granted_niosII_system_burst_5_upstream) OR cpu_data_master_granted_niosII_system_burst_6_upstream) OR cpu_data_master_granted_niosII_system_burst_7_upstream) OR cpu_data_master_granted_niosII_system_burst_8_upstream) OR cpu_data_master_granted_niosII_system_burst_9_upstream;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_cpu_data_master_readdatavalid <= (((((((((((((((cpu_data_master_read_data_valid_niosII_system_burst_1_upstream OR ((cpu_data_master_read_data_valid_niosII_system_burst_11_upstream AND dbs_rdv_counter_overflow))) OR ((cpu_data_master_read_data_valid_niosII_system_burst_13_upstream AND dbs_rdv_counter_overflow))) OR cpu_data_master_read_data_valid_niosII_system_burst_14_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_15_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_16_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_17_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_18_upstream) OR ((cpu_data_master_read_data_valid_niosII_system_burst_20_upstream AND dbs_rdv_counter_overflow))) OR cpu_data_master_read_data_valid_niosII_system_burst_21_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_3_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_4_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_5_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_6_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_7_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_8_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_9_upstream;
  --latent slave read data valid which is not flushed, which is an e_mux
  cpu_data_master_readdatavalid <= ((((((((((((((((((((((((((((((((cpu_data_master_read_but_no_slave_selected OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid;
  --cpu/data_master readdata mux, which is an e_mux
  cpu_data_master_readdata <= (((((((((((((((((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_1_upstream, 32) OR niosII_system_burst_1_upstream_readdata_from_sa)) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_11_upstream, 32) OR Std_Logic_Vector'(niosII_system_burst_11_upstream_readdata_from_sa(15 DOWNTO 0) & dbs_latent_16_reg_segment_0)))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_13_upstream, 32) OR Std_Logic_Vector'(niosII_system_burst_13_upstream_readdata_from_sa(7 DOWNTO 0) & dbs_latent_8_reg_segment_2 & dbs_latent_8_reg_segment_1 & dbs_latent_8_reg_segment_0)))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_14_upstream, 32) OR (std_logic_vector'("0000000000000000") & (niosII_system_burst_14_upstream_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_15_upstream, 32) OR (std_logic_vector'("0000000000000000") & (niosII_system_burst_15_upstream_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_16_upstream, 32) OR (std_logic_vector'("0000000000000000") & (niosII_system_burst_16_upstream_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_17_upstream, 32) OR (std_logic_vector'("0000000000000000") & (niosII_system_burst_17_upstream_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_18_upstream, 32) OR (std_logic_vector'("0000000000000000") & (niosII_system_burst_18_upstream_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_20_upstream, 32) OR Std_Logic_Vector'(niosII_system_burst_20_upstream_readdata_from_sa(15 DOWNTO 0) & dbs_latent_16_reg_segment_0)))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_21_upstream, 32) OR niosII_system_burst_21_upstream_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_3_upstream, 32) OR niosII_system_burst_3_upstream_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_4_upstream, 32) OR niosII_system_burst_4_upstream_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_5_upstream, 32) OR (std_logic_vector'("0000000000000000") & (niosII_system_burst_5_upstream_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_6_upstream, 32) OR niosII_system_burst_6_upstream_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_7_upstream, 32) OR (std_logic_vector'("000000000000000000000000") & (niosII_system_burst_7_upstream_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_8_upstream, 32) OR (std_logic_vector'("000000000000000000000000") & (niosII_system_burst_8_upstream_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_read_data_valid_niosII_system_burst_9_upstream, 32) OR (std_logic_vector'("000000000000000000000000") & (niosII_system_burst_9_upstream_readdata_from_sa))));
  --actual waitrequest port, which is an e_assign
  internal_cpu_data_master_waitrequest <= NOT cpu_data_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_data_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_cpu_data_master_latency_counter <= p1_cpu_data_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_cpu_data_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((cpu_data_master_run AND cpu_data_master_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_cpu_data_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --input to latent dbs-16 stored 0, which is an e_mux
  p1_dbs_latent_16_reg_segment_0 <= A_WE_StdLogicVector((std_logic'((cpu_data_master_read_data_valid_niosII_system_burst_11_upstream)) = '1'), niosII_system_burst_11_upstream_readdata_from_sa, niosII_system_burst_20_upstream_readdata_from_sa);
  --dbs register for latent dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_data_master_dbs_rdv_counter(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
      end if;
    end if;

  end process;

  --mux write dbs 1, which is an e_mux
  cpu_data_master_dbs_write_16 <= A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_dbs_address(1))) = '1'), cpu_data_master_writedata(31 DOWNTO 16), A_WE_StdLogicVector((std_logic'((NOT (internal_cpu_data_master_dbs_address(1)))) = '1'), cpu_data_master_writedata(15 DOWNTO 0), A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_dbs_address(1))) = '1'), cpu_data_master_writedata(31 DOWNTO 16), cpu_data_master_writedata(15 DOWNTO 0))));
  --dbs count increment, which is an e_mux
  cpu_data_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((cpu_data_master_requests_niosII_system_burst_11_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((cpu_data_master_requests_niosII_system_burst_13_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((cpu_data_master_requests_niosII_system_burst_20_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")))), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_cpu_data_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_cpu_data_master_dbs_address)) + (std_logic_vector'("0") & (cpu_data_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_data_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_cpu_data_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  cpu_data_master_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (cpu_data_master_dbs_rdv_counter)) + (std_logic_vector'("0") & (cpu_data_master_dbs_rdv_counter_inc))), 2);
  --cpu_data_master_rdv_inc_mux, which is an e_mux
  cpu_data_master_dbs_rdv_counter_inc <= A_EXT (A_WE_StdLogicVector((std_logic'((cpu_data_master_read_data_valid_niosII_system_burst_11_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((cpu_data_master_read_data_valid_niosII_system_burst_13_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000001"), std_logic_vector'("00000000000000000000000000000010"))), 2);
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream OR cpu_data_master_read_data_valid_niosII_system_burst_13_upstream) OR cpu_data_master_read_data_valid_niosII_system_burst_20_upstream;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_dbs_rdv_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        cpu_data_master_dbs_rdv_counter <= cpu_data_master_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= cpu_data_master_dbs_rdv_counter(1) AND NOT cpu_data_master_next_dbs_rdv_counter(1);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_data_master_granted_niosII_system_burst_11_upstream AND cpu_data_master_read)))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_11_upstream_waitrequest_from_sa))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_data_master_granted_niosII_system_burst_11_upstream AND cpu_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_11_upstream_waitrequest_from_sa)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_data_master_granted_niosII_system_burst_13_upstream AND cpu_data_master_read)))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_13_upstream_waitrequest_from_sa)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_data_master_granted_niosII_system_burst_13_upstream AND cpu_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_13_upstream_waitrequest_from_sa)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_data_master_granted_niosII_system_burst_20_upstream AND cpu_data_master_read)))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_20_upstream_waitrequest_from_sa)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_data_master_granted_niosII_system_burst_20_upstream AND cpu_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_20_upstream_waitrequest_from_sa)))))));
  --input to latent dbs-8 stored 0, which is an e_mux
  p1_dbs_latent_8_reg_segment_0 <= niosII_system_burst_13_upstream_readdata_from_sa;
  --dbs register for latent dbs-8 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_8_reg_segment_0 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((cpu_data_master_dbs_rdv_counter(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_8_reg_segment_0 <= p1_dbs_latent_8_reg_segment_0;
      end if;
    end if;

  end process;

  --input to latent dbs-8 stored 1, which is an e_mux
  p1_dbs_latent_8_reg_segment_1 <= niosII_system_burst_13_upstream_readdata_from_sa;
  --dbs register for latent dbs-8 segment 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_8_reg_segment_1 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((cpu_data_master_dbs_rdv_counter(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000001")))))) = '1' then 
        dbs_latent_8_reg_segment_1 <= p1_dbs_latent_8_reg_segment_1;
      end if;
    end if;

  end process;

  --input to latent dbs-8 stored 2, which is an e_mux
  p1_dbs_latent_8_reg_segment_2 <= niosII_system_burst_13_upstream_readdata_from_sa;
  --dbs register for latent dbs-8 segment 2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_8_reg_segment_2 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((cpu_data_master_dbs_rdv_counter(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000010")))))) = '1' then 
        dbs_latent_8_reg_segment_2 <= p1_dbs_latent_8_reg_segment_2;
      end if;
    end if;

  end process;

  --mux write dbs 2, which is an e_mux
  cpu_data_master_dbs_write_8 <= A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), cpu_data_master_writedata(7 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), cpu_data_master_writedata(15 DOWNTO 8), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), cpu_data_master_writedata(23 DOWNTO 16), cpu_data_master_writedata(31 DOWNTO 24))));
  --vhdl renameroo for output signals
  cpu_data_master_address_to_slave <= internal_cpu_data_master_address_to_slave;
  --vhdl renameroo for output signals
  cpu_data_master_dbs_address <= internal_cpu_data_master_dbs_address;
  --vhdl renameroo for output signals
  cpu_data_master_latency_counter <= internal_cpu_data_master_latency_counter;
  --vhdl renameroo for output signals
  cpu_data_master_waitrequest <= internal_cpu_data_master_waitrequest;
--synthesis translate_off
    --cpu_data_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_data_master_address_last_time <= cpu_data_master_address;
      end if;

    end process;

    --cpu/data_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpu_data_master_waitrequest AND ((cpu_data_master_read OR cpu_data_master_write));
      end if;

    end process;

    --cpu_data_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line6 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_data_master_address /= cpu_data_master_address_last_time))))) = '1' then 
          write(write_line6, now);
          write(write_line6, string'(": "));
          write(write_line6, string'("cpu_data_master_address did not heed wait!!!"));
          write(output, write_line6.all);
          deallocate (write_line6);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_data_master_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_burstcount_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        cpu_data_master_burstcount_last_time <= cpu_data_master_burstcount;
      end if;

    end process;

    --cpu_data_master_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line7 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_data_master_burstcount /= cpu_data_master_burstcount_last_time))))) = '1' then 
          write(write_line7, now);
          write(write_line7, string'(": "));
          write(write_line7, string'("cpu_data_master_burstcount did not heed wait!!!"));
          write(output, write_line7.all);
          deallocate (write_line7);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_data_master_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        cpu_data_master_byteenable_last_time <= cpu_data_master_byteenable;
      end if;

    end process;

    --cpu_data_master_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line8 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_data_master_byteenable /= cpu_data_master_byteenable_last_time))))) = '1' then 
          write(write_line8, now);
          write(write_line8, string'(": "));
          write(write_line8, string'("cpu_data_master_byteenable did not heed wait!!!"));
          write(output, write_line8.all);
          deallocate (write_line8);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_data_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_data_master_read_last_time <= cpu_data_master_read;
      end if;

    end process;

    --cpu_data_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line9 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_data_master_read) /= std_logic'(cpu_data_master_read_last_time)))))) = '1' then 
          write(write_line9, now);
          write(write_line9, string'(": "));
          write(write_line9, string'("cpu_data_master_read did not heed wait!!!"));
          write(output, write_line9.all);
          deallocate (write_line9);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_data_master_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_data_master_write_last_time <= cpu_data_master_write;
      end if;

    end process;

    --cpu_data_master_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line10 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_data_master_write) /= std_logic'(cpu_data_master_write_last_time)))))) = '1' then 
          write(write_line10, now);
          write(write_line10, string'(": "));
          write(write_line10, string'("cpu_data_master_write did not heed wait!!!"));
          write(output, write_line10.all);
          deallocate (write_line10);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_data_master_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_data_master_writedata_last_time <= cpu_data_master_writedata;
      end if;

    end process;

    --cpu_data_master_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line11 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((cpu_data_master_writedata /= cpu_data_master_writedata_last_time)))) AND cpu_data_master_write)) = '1' then 
          write(write_line11, now);
          write(write_line11, string'(": "));
          write(write_line11, string'("cpu_data_master_writedata did not heed wait!!!"));
          write(output, write_line11.all);
          deallocate (write_line11);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_instruction_master_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_instruction_master_granted_niosII_system_burst_0_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_granted_niosII_system_burst_10_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_granted_niosII_system_burst_12_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_granted_niosII_system_burst_19_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_granted_niosII_system_burst_2_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_requests_niosII_system_burst_0_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_requests_niosII_system_burst_10_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_requests_niosII_system_burst_12_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_requests_niosII_system_burst_19_upstream : IN STD_LOGIC;
                 signal cpu_instruction_master_requests_niosII_system_burst_2_upstream : IN STD_LOGIC;
                 signal d1_niosII_system_burst_0_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_10_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_12_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_19_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_system_burst_2_upstream_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_0_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_0_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_10_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_10_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_12_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_12_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_19_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_19_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_2_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_2_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : OUT STD_LOGIC;
                 signal cpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                 signal cpu_instruction_master_waitrequest : OUT STD_LOGIC
              );
end entity cpu_instruction_master_arbitrator;


architecture europa of cpu_instruction_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpu_instruction_master_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_instruction_master_burstcount_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_instruction_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_is_granted_some_slave :  STD_LOGIC;
                signal cpu_instruction_master_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_read_but_no_slave_selected :  STD_LOGIC;
                signal cpu_instruction_master_read_last_time :  STD_LOGIC;
                signal cpu_instruction_master_run :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_latent_8_reg_segment_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_latent_8_reg_segment_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_latent_8_reg_segment_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_cpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_cpu_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_instruction_master_latency_counter :  STD_LOGIC;
                signal internal_cpu_instruction_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_cpu_instruction_master_latency_counter :  STD_LOGIC;
                signal p1_dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_dbs_latent_8_reg_segment_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_dbs_latent_8_reg_segment_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_dbs_latent_8_reg_segment_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_cpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream OR NOT cpu_instruction_master_requests_niosII_system_burst_0_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream OR NOT (cpu_instruction_master_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_0_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_read))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream OR NOT cpu_instruction_master_requests_niosII_system_burst_10_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream OR NOT cpu_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_10_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_read)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream OR NOT cpu_instruction_master_requests_niosII_system_burst_12_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream OR NOT cpu_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_12_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_read)))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_instruction_master_run <= r_0 AND r_1;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream OR NOT cpu_instruction_master_requests_niosII_system_burst_19_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream OR NOT cpu_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_19_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_read)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream OR NOT cpu_instruction_master_requests_niosII_system_burst_2_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream OR NOT (cpu_instruction_master_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_2_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_read))))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_instruction_master_address_to_slave <= cpu_instruction_master_address(24 DOWNTO 0);
  --cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_instruction_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_instruction_master_read_but_no_slave_selected <= (cpu_instruction_master_read AND cpu_instruction_master_run) AND NOT cpu_instruction_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  cpu_instruction_master_is_granted_some_slave <= (((cpu_instruction_master_granted_niosII_system_burst_0_upstream OR cpu_instruction_master_granted_niosII_system_burst_10_upstream) OR cpu_instruction_master_granted_niosII_system_burst_12_upstream) OR cpu_instruction_master_granted_niosII_system_burst_19_upstream) OR cpu_instruction_master_granted_niosII_system_burst_2_upstream;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_cpu_instruction_master_readdatavalid <= (((cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream OR ((cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream AND dbs_rdv_counter_overflow))) OR ((cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream AND dbs_rdv_counter_overflow))) OR ((cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream AND dbs_rdv_counter_overflow))) OR cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream;
  --latent slave read data valid which is not flushed, which is an e_mux
  cpu_instruction_master_readdatavalid <= ((((((((cpu_instruction_master_read_but_no_slave_selected OR pre_flush_cpu_instruction_master_readdatavalid) OR cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_cpu_instruction_master_readdatavalid) OR cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_cpu_instruction_master_readdatavalid) OR cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_cpu_instruction_master_readdatavalid) OR cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_cpu_instruction_master_readdatavalid;
  --cpu/instruction_master readdata mux, which is an e_mux
  cpu_instruction_master_readdata <= (((((A_REP(NOT cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream, 32) OR niosII_system_burst_0_upstream_readdata_from_sa)) AND ((A_REP(NOT cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream, 32) OR Std_Logic_Vector'(niosII_system_burst_10_upstream_readdata_from_sa(15 DOWNTO 0) & dbs_latent_16_reg_segment_0)))) AND ((A_REP(NOT cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream, 32) OR Std_Logic_Vector'(niosII_system_burst_12_upstream_readdata_from_sa(7 DOWNTO 0) & dbs_latent_8_reg_segment_2 & dbs_latent_8_reg_segment_1 & dbs_latent_8_reg_segment_0)))) AND ((A_REP(NOT cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream, 32) OR Std_Logic_Vector'(niosII_system_burst_19_upstream_readdata_from_sa(15 DOWNTO 0) & dbs_latent_16_reg_segment_0)))) AND ((A_REP(NOT cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream, 32) OR niosII_system_burst_2_upstream_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_cpu_instruction_master_waitrequest <= NOT cpu_instruction_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_instruction_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_cpu_instruction_master_latency_counter <= p1_cpu_instruction_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_cpu_instruction_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((cpu_instruction_master_run AND cpu_instruction_master_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_cpu_instruction_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --input to latent dbs-16 stored 0, which is an e_mux
  p1_dbs_latent_16_reg_segment_0 <= A_WE_StdLogicVector((std_logic'((cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream)) = '1'), niosII_system_burst_10_upstream_readdata_from_sa, niosII_system_burst_19_upstream_readdata_from_sa);
  --dbs register for latent dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_dbs_rdv_counter(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
      end if;
    end if;

  end process;

  --dbs count increment, which is an e_mux
  cpu_instruction_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((cpu_instruction_master_requests_niosII_system_burst_10_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((cpu_instruction_master_requests_niosII_system_burst_12_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((cpu_instruction_master_requests_niosII_system_burst_19_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")))), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_cpu_instruction_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_cpu_instruction_master_dbs_address)) + (std_logic_vector'("0") & (cpu_instruction_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_instruction_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_cpu_instruction_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  cpu_instruction_master_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (cpu_instruction_master_dbs_rdv_counter)) + (std_logic_vector'("0") & (cpu_instruction_master_dbs_rdv_counter_inc))), 2);
  --cpu_instruction_master_rdv_inc_mux, which is an e_mux
  cpu_instruction_master_dbs_rdv_counter_inc <= A_EXT (A_WE_StdLogicVector((std_logic'((cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000001"), std_logic_vector'("00000000000000000000000000000010"))), 2);
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= (cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream OR cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream) OR cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_instruction_master_dbs_rdv_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        cpu_instruction_master_dbs_rdv_counter <= cpu_instruction_master_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= cpu_instruction_master_dbs_rdv_counter(1) AND NOT cpu_instruction_master_next_dbs_rdv_counter(1);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_granted_niosII_system_burst_10_upstream AND cpu_instruction_master_read)))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_10_upstream_waitrequest_from_sa))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_granted_niosII_system_burst_12_upstream AND cpu_instruction_master_read)))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_12_upstream_waitrequest_from_sa)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_granted_niosII_system_burst_19_upstream AND cpu_instruction_master_read)))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_19_upstream_waitrequest_from_sa)))))));
  --input to latent dbs-8 stored 0, which is an e_mux
  p1_dbs_latent_8_reg_segment_0 <= niosII_system_burst_12_upstream_readdata_from_sa;
  --dbs register for latent dbs-8 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_8_reg_segment_0 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((cpu_instruction_master_dbs_rdv_counter(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_8_reg_segment_0 <= p1_dbs_latent_8_reg_segment_0;
      end if;
    end if;

  end process;

  --input to latent dbs-8 stored 1, which is an e_mux
  p1_dbs_latent_8_reg_segment_1 <= niosII_system_burst_12_upstream_readdata_from_sa;
  --dbs register for latent dbs-8 segment 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_8_reg_segment_1 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((cpu_instruction_master_dbs_rdv_counter(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000001")))))) = '1' then 
        dbs_latent_8_reg_segment_1 <= p1_dbs_latent_8_reg_segment_1;
      end if;
    end if;

  end process;

  --input to latent dbs-8 stored 2, which is an e_mux
  p1_dbs_latent_8_reg_segment_2 <= niosII_system_burst_12_upstream_readdata_from_sa;
  --dbs register for latent dbs-8 segment 2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_8_reg_segment_2 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((cpu_instruction_master_dbs_rdv_counter(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000010")))))) = '1' then 
        dbs_latent_8_reg_segment_2 <= p1_dbs_latent_8_reg_segment_2;
      end if;
    end if;

  end process;

  --vhdl renameroo for output signals
  cpu_instruction_master_address_to_slave <= internal_cpu_instruction_master_address_to_slave;
  --vhdl renameroo for output signals
  cpu_instruction_master_dbs_address <= internal_cpu_instruction_master_dbs_address;
  --vhdl renameroo for output signals
  cpu_instruction_master_latency_counter <= internal_cpu_instruction_master_latency_counter;
  --vhdl renameroo for output signals
  cpu_instruction_master_waitrequest <= internal_cpu_instruction_master_waitrequest;
--synthesis translate_off
    --cpu_instruction_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_instruction_master_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_instruction_master_address_last_time <= cpu_instruction_master_address;
      end if;

    end process;

    --cpu/instruction_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpu_instruction_master_waitrequest AND (cpu_instruction_master_read);
      end if;

    end process;

    --cpu_instruction_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line12 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_instruction_master_address /= cpu_instruction_master_address_last_time))))) = '1' then 
          write(write_line12, now);
          write(write_line12, string'(": "));
          write(write_line12, string'("cpu_instruction_master_address did not heed wait!!!"));
          write(output, write_line12.all);
          deallocate (write_line12);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_instruction_master_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_instruction_master_burstcount_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        cpu_instruction_master_burstcount_last_time <= cpu_instruction_master_burstcount;
      end if;

    end process;

    --cpu_instruction_master_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line13 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_instruction_master_burstcount /= cpu_instruction_master_burstcount_last_time))))) = '1' then 
          write(write_line13, now);
          write(write_line13, string'(": "));
          write(write_line13, string'("cpu_instruction_master_burstcount did not heed wait!!!"));
          write(output, write_line13.all);
          deallocate (write_line13);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_instruction_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_instruction_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_instruction_master_read_last_time <= cpu_instruction_master_read;
      end if;

    end process;

    --cpu_instruction_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line14 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_instruction_master_read) /= std_logic'(cpu_instruction_master_read_last_time)))))) = '1' then 
          write(write_line14, now);
          write(write_line14, string'(": "));
          write(write_line14, string'("cpu_instruction_master_read did not heed wait!!!"));
          write(output, write_line14.all);
          deallocate (write_line14);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity dm9000a_inst_avalon_slave_0_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_irq : IN STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_16_downstream_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_16_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_16_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_16_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_dm9000a_inst_avalon_slave_0_end_xfer : OUT STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_address : OUT STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_chipselect_n : OUT STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_irq_from_sa : OUT STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_read_n : OUT STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal dm9000a_inst_avalon_slave_0_reset_n : OUT STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_write_n : OUT STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 : OUT STD_LOGIC;
                 signal niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 : OUT STD_LOGIC;
                 signal niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0 : OUT STD_LOGIC;
                 signal niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 : OUT STD_LOGIC
              );
end entity dm9000a_inst_avalon_slave_0_arbitrator;


architecture europa of dm9000a_inst_avalon_slave_0_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_allgrants :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_allow_new_arb_cycle :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_any_bursting_master_saved_grant :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_any_continuerequest :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_arb_counter_enable :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_arb_share_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal dm9000a_inst_avalon_slave_0_arb_share_counter_next_value :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal dm9000a_inst_avalon_slave_0_arb_share_set_values :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal dm9000a_inst_avalon_slave_0_beginbursttransfer_internal :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_begins_xfer :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_end_xfer :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_firsttransfer :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_grant_vector :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_in_a_read_cycle :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_in_a_write_cycle :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_master_qreq_vector :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_non_bursting_master_requests :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_reg_firsttransfer :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_slavearbiterlockenable :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_slavearbiterlockenable2 :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_unreg_firsttransfer :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_waits_for_read :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_waits_for_write :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_dm9000a_inst_avalon_slave_0 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 :  STD_LOGIC;
                signal internal_niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 :  STD_LOGIC;
                signal internal_niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_saved_grant_dm9000a_inst_avalon_slave_0 :  STD_LOGIC;
                signal wait_for_dm9000a_inst_avalon_slave_0_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT dm9000a_inst_avalon_slave_0_end_xfer;
    end if;

  end process;

  dm9000a_inst_avalon_slave_0_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0);
  --assign dm9000a_inst_avalon_slave_0_readdata_from_sa = dm9000a_inst_avalon_slave_0_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  dm9000a_inst_avalon_slave_0_readdata_from_sa <= dm9000a_inst_avalon_slave_0_readdata;
  internal_niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_16_downstream_read OR niosII_system_burst_16_downstream_write)))))));
  --dm9000a_inst_avalon_slave_0_arb_share_counter set values, which is an e_mux
  dm9000a_inst_avalon_slave_0_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_16_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --dm9000a_inst_avalon_slave_0_non_bursting_master_requests mux, which is an e_mux
  dm9000a_inst_avalon_slave_0_non_bursting_master_requests <= std_logic'('0');
  --dm9000a_inst_avalon_slave_0_any_bursting_master_saved_grant mux, which is an e_mux
  dm9000a_inst_avalon_slave_0_any_bursting_master_saved_grant <= niosII_system_burst_16_downstream_saved_grant_dm9000a_inst_avalon_slave_0;
  --dm9000a_inst_avalon_slave_0_arb_share_counter_next_value assignment, which is an e_assign
  dm9000a_inst_avalon_slave_0_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(dm9000a_inst_avalon_slave_0_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (dm9000a_inst_avalon_slave_0_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(dm9000a_inst_avalon_slave_0_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (dm9000a_inst_avalon_slave_0_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 5);
  --dm9000a_inst_avalon_slave_0_allgrants all slave grants, which is an e_mux
  dm9000a_inst_avalon_slave_0_allgrants <= dm9000a_inst_avalon_slave_0_grant_vector;
  --dm9000a_inst_avalon_slave_0_end_xfer assignment, which is an e_assign
  dm9000a_inst_avalon_slave_0_end_xfer <= NOT ((dm9000a_inst_avalon_slave_0_waits_for_read OR dm9000a_inst_avalon_slave_0_waits_for_write));
  --end_xfer_arb_share_counter_term_dm9000a_inst_avalon_slave_0 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_dm9000a_inst_avalon_slave_0 <= dm9000a_inst_avalon_slave_0_end_xfer AND (((NOT dm9000a_inst_avalon_slave_0_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --dm9000a_inst_avalon_slave_0_arb_share_counter arbitration counter enable, which is an e_assign
  dm9000a_inst_avalon_slave_0_arb_counter_enable <= ((end_xfer_arb_share_counter_term_dm9000a_inst_avalon_slave_0 AND dm9000a_inst_avalon_slave_0_allgrants)) OR ((end_xfer_arb_share_counter_term_dm9000a_inst_avalon_slave_0 AND NOT dm9000a_inst_avalon_slave_0_non_bursting_master_requests));
  --dm9000a_inst_avalon_slave_0_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dm9000a_inst_avalon_slave_0_arb_share_counter <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(dm9000a_inst_avalon_slave_0_arb_counter_enable) = '1' then 
        dm9000a_inst_avalon_slave_0_arb_share_counter <= dm9000a_inst_avalon_slave_0_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --dm9000a_inst_avalon_slave_0_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dm9000a_inst_avalon_slave_0_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((dm9000a_inst_avalon_slave_0_master_qreq_vector AND end_xfer_arb_share_counter_term_dm9000a_inst_avalon_slave_0)) OR ((end_xfer_arb_share_counter_term_dm9000a_inst_avalon_slave_0 AND NOT dm9000a_inst_avalon_slave_0_non_bursting_master_requests)))) = '1' then 
        dm9000a_inst_avalon_slave_0_slavearbiterlockenable <= or_reduce(dm9000a_inst_avalon_slave_0_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_16/downstream dm9000a_inst/avalon_slave_0 arbiterlock, which is an e_assign
  niosII_system_burst_16_downstream_arbiterlock <= dm9000a_inst_avalon_slave_0_slavearbiterlockenable AND niosII_system_burst_16_downstream_continuerequest;
  --dm9000a_inst_avalon_slave_0_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  dm9000a_inst_avalon_slave_0_slavearbiterlockenable2 <= or_reduce(dm9000a_inst_avalon_slave_0_arb_share_counter_next_value);
  --niosII_system_burst_16/downstream dm9000a_inst/avalon_slave_0 arbiterlock2, which is an e_assign
  niosII_system_burst_16_downstream_arbiterlock2 <= dm9000a_inst_avalon_slave_0_slavearbiterlockenable2 AND niosII_system_burst_16_downstream_continuerequest;
  --dm9000a_inst_avalon_slave_0_any_continuerequest at least one master continues requesting, which is an e_assign
  dm9000a_inst_avalon_slave_0_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_16_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_16_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 <= internal_niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 AND NOT ((niosII_system_burst_16_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_16_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0, which is an e_mux
  niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0 <= (internal_niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 AND niosII_system_burst_16_downstream_read) AND NOT dm9000a_inst_avalon_slave_0_waits_for_read;
  --dm9000a_inst_avalon_slave_0_writedata mux, which is an e_mux
  dm9000a_inst_avalon_slave_0_writedata <= niosII_system_burst_16_downstream_writedata;
  --master is always granted when requested
  internal_niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 <= internal_niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0;
  --niosII_system_burst_16/downstream saved-grant dm9000a_inst/avalon_slave_0, which is an e_assign
  niosII_system_burst_16_downstream_saved_grant_dm9000a_inst_avalon_slave_0 <= internal_niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0;
  --allow new arb cycle for dm9000a_inst/avalon_slave_0, which is an e_assign
  dm9000a_inst_avalon_slave_0_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  dm9000a_inst_avalon_slave_0_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  dm9000a_inst_avalon_slave_0_master_qreq_vector <= std_logic'('1');
  --dm9000a_inst_avalon_slave_0_reset_n assignment, which is an e_assign
  dm9000a_inst_avalon_slave_0_reset_n <= reset_n;
  dm9000a_inst_avalon_slave_0_chipselect_n <= NOT internal_niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0;
  --dm9000a_inst_avalon_slave_0_firsttransfer first transaction, which is an e_assign
  dm9000a_inst_avalon_slave_0_firsttransfer <= A_WE_StdLogic((std_logic'(dm9000a_inst_avalon_slave_0_begins_xfer) = '1'), dm9000a_inst_avalon_slave_0_unreg_firsttransfer, dm9000a_inst_avalon_slave_0_reg_firsttransfer);
  --dm9000a_inst_avalon_slave_0_unreg_firsttransfer first transaction, which is an e_assign
  dm9000a_inst_avalon_slave_0_unreg_firsttransfer <= NOT ((dm9000a_inst_avalon_slave_0_slavearbiterlockenable AND dm9000a_inst_avalon_slave_0_any_continuerequest));
  --dm9000a_inst_avalon_slave_0_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dm9000a_inst_avalon_slave_0_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(dm9000a_inst_avalon_slave_0_begins_xfer) = '1' then 
        dm9000a_inst_avalon_slave_0_reg_firsttransfer <= dm9000a_inst_avalon_slave_0_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --dm9000a_inst_avalon_slave_0_beginbursttransfer_internal begin burst transfer, which is an e_assign
  dm9000a_inst_avalon_slave_0_beginbursttransfer_internal <= dm9000a_inst_avalon_slave_0_begins_xfer;
  --~dm9000a_inst_avalon_slave_0_read_n assignment, which is an e_mux
  dm9000a_inst_avalon_slave_0_read_n <= NOT ((internal_niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 AND niosII_system_burst_16_downstream_read));
  --~dm9000a_inst_avalon_slave_0_write_n assignment, which is an e_mux
  dm9000a_inst_avalon_slave_0_write_n <= NOT ((internal_niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 AND niosII_system_burst_16_downstream_write));
  --dm9000a_inst_avalon_slave_0_address mux, which is an e_mux
  dm9000a_inst_avalon_slave_0_address <= niosII_system_burst_16_downstream_nativeaddress(0);
  --d1_dm9000a_inst_avalon_slave_0_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_dm9000a_inst_avalon_slave_0_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_dm9000a_inst_avalon_slave_0_end_xfer <= dm9000a_inst_avalon_slave_0_end_xfer;
    end if;

  end process;

  --dm9000a_inst_avalon_slave_0_waits_for_read in a cycle, which is an e_mux
  dm9000a_inst_avalon_slave_0_waits_for_read <= dm9000a_inst_avalon_slave_0_in_a_read_cycle AND dm9000a_inst_avalon_slave_0_begins_xfer;
  --dm9000a_inst_avalon_slave_0_in_a_read_cycle assignment, which is an e_assign
  dm9000a_inst_avalon_slave_0_in_a_read_cycle <= internal_niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 AND niosII_system_burst_16_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= dm9000a_inst_avalon_slave_0_in_a_read_cycle;
  --dm9000a_inst_avalon_slave_0_waits_for_write in a cycle, which is an e_mux
  dm9000a_inst_avalon_slave_0_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dm9000a_inst_avalon_slave_0_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --dm9000a_inst_avalon_slave_0_in_a_write_cycle assignment, which is an e_assign
  dm9000a_inst_avalon_slave_0_in_a_write_cycle <= internal_niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 AND niosII_system_burst_16_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= dm9000a_inst_avalon_slave_0_in_a_write_cycle;
  wait_for_dm9000a_inst_avalon_slave_0_counter <= std_logic'('0');
  --assign dm9000a_inst_avalon_slave_0_irq_from_sa = dm9000a_inst_avalon_slave_0_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  dm9000a_inst_avalon_slave_0_irq_from_sa <= dm9000a_inst_avalon_slave_0_irq;
  --vhdl renameroo for output signals
  niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 <= internal_niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0;
  --vhdl renameroo for output signals
  niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 <= internal_niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0;
  --vhdl renameroo for output signals
  niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 <= internal_niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0;
--synthesis translate_off
    --dm9000a_inst/avalon_slave_0 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_16/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line15 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_16_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line15, now);
          write(write_line15, string'(": "));
          write(write_line15, string'("niosII_system_burst_16/downstream drove 0 on its 'arbitrationshare' port while accessing slave dm9000a_inst/avalon_slave_0"));
          write(output, write_line15.all);
          deallocate (write_line15);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_16/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line16 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_16_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line16, now);
          write(write_line16, string'(": "));
          write(write_line16, string'("niosII_system_burst_16/downstream drove 0 on its 'burstcount' port while accessing slave dm9000a_inst/avalon_slave_0"));
          write(output, write_line16.all);
          deallocate (write_line16);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity high_res_timer_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal high_res_timer_s1_irq : IN STD_LOGIC;
                 signal high_res_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_15_downstream_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_15_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_15_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_15_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_high_res_timer_s1_end_xfer : OUT STD_LOGIC;
                 signal high_res_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal high_res_timer_s1_chipselect : OUT STD_LOGIC;
                 signal high_res_timer_s1_irq_from_sa : OUT STD_LOGIC;
                 signal high_res_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal high_res_timer_s1_reset_n : OUT STD_LOGIC;
                 signal high_res_timer_s1_write_n : OUT STD_LOGIC;
                 signal high_res_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_15_downstream_granted_high_res_timer_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_15_downstream_requests_high_res_timer_s1 : OUT STD_LOGIC
              );
end entity high_res_timer_s1_arbitrator;


architecture europa of high_res_timer_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_high_res_timer_s1 :  STD_LOGIC;
                signal high_res_timer_s1_allgrants :  STD_LOGIC;
                signal high_res_timer_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal high_res_timer_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal high_res_timer_s1_any_continuerequest :  STD_LOGIC;
                signal high_res_timer_s1_arb_counter_enable :  STD_LOGIC;
                signal high_res_timer_s1_arb_share_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal high_res_timer_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal high_res_timer_s1_arb_share_set_values :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal high_res_timer_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal high_res_timer_s1_begins_xfer :  STD_LOGIC;
                signal high_res_timer_s1_end_xfer :  STD_LOGIC;
                signal high_res_timer_s1_firsttransfer :  STD_LOGIC;
                signal high_res_timer_s1_grant_vector :  STD_LOGIC;
                signal high_res_timer_s1_in_a_read_cycle :  STD_LOGIC;
                signal high_res_timer_s1_in_a_write_cycle :  STD_LOGIC;
                signal high_res_timer_s1_master_qreq_vector :  STD_LOGIC;
                signal high_res_timer_s1_non_bursting_master_requests :  STD_LOGIC;
                signal high_res_timer_s1_reg_firsttransfer :  STD_LOGIC;
                signal high_res_timer_s1_slavearbiterlockenable :  STD_LOGIC;
                signal high_res_timer_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal high_res_timer_s1_unreg_firsttransfer :  STD_LOGIC;
                signal high_res_timer_s1_waits_for_read :  STD_LOGIC;
                signal high_res_timer_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_15_downstream_granted_high_res_timer_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_15_downstream_requests_high_res_timer_s1 :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_saved_grant_high_res_timer_s1 :  STD_LOGIC;
                signal wait_for_high_res_timer_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT high_res_timer_s1_end_xfer;
    end if;

  end process;

  high_res_timer_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1);
  --assign high_res_timer_s1_readdata_from_sa = high_res_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  high_res_timer_s1_readdata_from_sa <= high_res_timer_s1_readdata;
  internal_niosII_system_burst_15_downstream_requests_high_res_timer_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_15_downstream_read OR niosII_system_burst_15_downstream_write)))))));
  --high_res_timer_s1_arb_share_counter set values, which is an e_mux
  high_res_timer_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_15_downstream_granted_high_res_timer_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_15_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --high_res_timer_s1_non_bursting_master_requests mux, which is an e_mux
  high_res_timer_s1_non_bursting_master_requests <= std_logic'('0');
  --high_res_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  high_res_timer_s1_any_bursting_master_saved_grant <= niosII_system_burst_15_downstream_saved_grant_high_res_timer_s1;
  --high_res_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  high_res_timer_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(high_res_timer_s1_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (high_res_timer_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(high_res_timer_s1_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (high_res_timer_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 5);
  --high_res_timer_s1_allgrants all slave grants, which is an e_mux
  high_res_timer_s1_allgrants <= high_res_timer_s1_grant_vector;
  --high_res_timer_s1_end_xfer assignment, which is an e_assign
  high_res_timer_s1_end_xfer <= NOT ((high_res_timer_s1_waits_for_read OR high_res_timer_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_high_res_timer_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_high_res_timer_s1 <= high_res_timer_s1_end_xfer AND (((NOT high_res_timer_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --high_res_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  high_res_timer_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_high_res_timer_s1 AND high_res_timer_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_high_res_timer_s1 AND NOT high_res_timer_s1_non_bursting_master_requests));
  --high_res_timer_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      high_res_timer_s1_arb_share_counter <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(high_res_timer_s1_arb_counter_enable) = '1' then 
        high_res_timer_s1_arb_share_counter <= high_res_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --high_res_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      high_res_timer_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((high_res_timer_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_high_res_timer_s1)) OR ((end_xfer_arb_share_counter_term_high_res_timer_s1 AND NOT high_res_timer_s1_non_bursting_master_requests)))) = '1' then 
        high_res_timer_s1_slavearbiterlockenable <= or_reduce(high_res_timer_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_15/downstream high_res_timer/s1 arbiterlock, which is an e_assign
  niosII_system_burst_15_downstream_arbiterlock <= high_res_timer_s1_slavearbiterlockenable AND niosII_system_burst_15_downstream_continuerequest;
  --high_res_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  high_res_timer_s1_slavearbiterlockenable2 <= or_reduce(high_res_timer_s1_arb_share_counter_next_value);
  --niosII_system_burst_15/downstream high_res_timer/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_15_downstream_arbiterlock2 <= high_res_timer_s1_slavearbiterlockenable2 AND niosII_system_burst_15_downstream_continuerequest;
  --high_res_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  high_res_timer_s1_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_15_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_15_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 <= internal_niosII_system_burst_15_downstream_requests_high_res_timer_s1 AND NOT ((niosII_system_burst_15_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_15_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1, which is an e_mux
  niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1 <= (internal_niosII_system_burst_15_downstream_granted_high_res_timer_s1 AND niosII_system_burst_15_downstream_read) AND NOT high_res_timer_s1_waits_for_read;
  --high_res_timer_s1_writedata mux, which is an e_mux
  high_res_timer_s1_writedata <= niosII_system_burst_15_downstream_writedata;
  --master is always granted when requested
  internal_niosII_system_burst_15_downstream_granted_high_res_timer_s1 <= internal_niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1;
  --niosII_system_burst_15/downstream saved-grant high_res_timer/s1, which is an e_assign
  niosII_system_burst_15_downstream_saved_grant_high_res_timer_s1 <= internal_niosII_system_burst_15_downstream_requests_high_res_timer_s1;
  --allow new arb cycle for high_res_timer/s1, which is an e_assign
  high_res_timer_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  high_res_timer_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  high_res_timer_s1_master_qreq_vector <= std_logic'('1');
  --high_res_timer_s1_reset_n assignment, which is an e_assign
  high_res_timer_s1_reset_n <= reset_n;
  high_res_timer_s1_chipselect <= internal_niosII_system_burst_15_downstream_granted_high_res_timer_s1;
  --high_res_timer_s1_firsttransfer first transaction, which is an e_assign
  high_res_timer_s1_firsttransfer <= A_WE_StdLogic((std_logic'(high_res_timer_s1_begins_xfer) = '1'), high_res_timer_s1_unreg_firsttransfer, high_res_timer_s1_reg_firsttransfer);
  --high_res_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  high_res_timer_s1_unreg_firsttransfer <= NOT ((high_res_timer_s1_slavearbiterlockenable AND high_res_timer_s1_any_continuerequest));
  --high_res_timer_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      high_res_timer_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(high_res_timer_s1_begins_xfer) = '1' then 
        high_res_timer_s1_reg_firsttransfer <= high_res_timer_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --high_res_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  high_res_timer_s1_beginbursttransfer_internal <= high_res_timer_s1_begins_xfer;
  --~high_res_timer_s1_write_n assignment, which is an e_mux
  high_res_timer_s1_write_n <= NOT ((internal_niosII_system_burst_15_downstream_granted_high_res_timer_s1 AND niosII_system_burst_15_downstream_write));
  --high_res_timer_s1_address mux, which is an e_mux
  high_res_timer_s1_address <= niosII_system_burst_15_downstream_nativeaddress (2 DOWNTO 0);
  --d1_high_res_timer_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_high_res_timer_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_high_res_timer_s1_end_xfer <= high_res_timer_s1_end_xfer;
    end if;

  end process;

  --high_res_timer_s1_waits_for_read in a cycle, which is an e_mux
  high_res_timer_s1_waits_for_read <= high_res_timer_s1_in_a_read_cycle AND high_res_timer_s1_begins_xfer;
  --high_res_timer_s1_in_a_read_cycle assignment, which is an e_assign
  high_res_timer_s1_in_a_read_cycle <= internal_niosII_system_burst_15_downstream_granted_high_res_timer_s1 AND niosII_system_burst_15_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= high_res_timer_s1_in_a_read_cycle;
  --high_res_timer_s1_waits_for_write in a cycle, which is an e_mux
  high_res_timer_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(high_res_timer_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --high_res_timer_s1_in_a_write_cycle assignment, which is an e_assign
  high_res_timer_s1_in_a_write_cycle <= internal_niosII_system_burst_15_downstream_granted_high_res_timer_s1 AND niosII_system_burst_15_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= high_res_timer_s1_in_a_write_cycle;
  wait_for_high_res_timer_s1_counter <= std_logic'('0');
  --assign high_res_timer_s1_irq_from_sa = high_res_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  high_res_timer_s1_irq_from_sa <= high_res_timer_s1_irq;
  --vhdl renameroo for output signals
  niosII_system_burst_15_downstream_granted_high_res_timer_s1 <= internal_niosII_system_burst_15_downstream_granted_high_res_timer_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 <= internal_niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_15_downstream_requests_high_res_timer_s1 <= internal_niosII_system_burst_15_downstream_requests_high_res_timer_s1;
--synthesis translate_off
    --high_res_timer/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_15/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line17 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_15_downstream_requests_high_res_timer_s1 AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_15_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line17, now);
          write(write_line17, string'(": "));
          write(write_line17, string'("niosII_system_burst_15/downstream drove 0 on its 'arbitrationshare' port while accessing slave high_res_timer/s1"));
          write(output, write_line17.all);
          deallocate (write_line17);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_15/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line18 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_15_downstream_requests_high_res_timer_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_15_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line18, now);
          write(write_line18, string'(": "));
          write(write_line18, string'("niosII_system_burst_15/downstream drove 0 on its 'burstcount' port while accessing slave high_res_timer/s1"));
          write(output, write_line18.all);
          deallocate (write_line18);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity jtag_uart_avalon_jtag_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_6_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_6_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_6_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC
              );
end entity jtag_uart_avalon_jtag_slave_arbitrator;


architecture europa of jtag_uart_avalon_jtag_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allgrants :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_continuerequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_counter_enable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_begins_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_grant_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_read_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_write_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_master_qreq_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_non_bursting_master_requests :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_unreg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_read :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_write :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_saved_grant_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal wait_for_jtag_uart_avalon_jtag_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  jtag_uart_avalon_jtag_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave);
  --assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readdata_from_sa <= jtag_uart_avalon_jtag_slave_readdata;
  internal_niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_6_downstream_read OR niosII_system_burst_6_downstream_write)))))));
  --assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_dataavailable_from_sa <= jtag_uart_avalon_jtag_slave_dataavailable;
  --assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readyfordata_from_sa <= jtag_uart_avalon_jtag_slave_readyfordata;
  --assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= jtag_uart_avalon_jtag_slave_waitrequest;
  --jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  jtag_uart_avalon_jtag_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_6_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_non_bursting_master_requests <= std_logic'('0');
  --jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant <= niosII_system_burst_6_downstream_saved_grant_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(jtag_uart_avalon_jtag_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (jtag_uart_avalon_jtag_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(jtag_uart_avalon_jtag_slave_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (jtag_uart_avalon_jtag_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  jtag_uart_avalon_jtag_slave_allgrants <= jtag_uart_avalon_jtag_slave_grant_vector;
  --jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_end_xfer <= NOT ((jtag_uart_avalon_jtag_slave_waits_for_read OR jtag_uart_avalon_jtag_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave <= jtag_uart_avalon_jtag_slave_end_xfer AND (((NOT jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND jtag_uart_avalon_jtag_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests));
  --jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_arb_counter_enable) = '1' then 
        jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((jtag_uart_avalon_jtag_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests)))) = '1' then 
        jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= or_reduce(jtag_uart_avalon_jtag_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_6/downstream jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  niosII_system_burst_6_downstream_arbiterlock <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND niosII_system_burst_6_downstream_continuerequest;
  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 <= or_reduce(jtag_uart_avalon_jtag_slave_arb_share_counter_next_value);
  --niosII_system_burst_6/downstream jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  niosII_system_burst_6_downstream_arbiterlock2 <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 AND niosII_system_burst_6_downstream_continuerequest;
  --jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  jtag_uart_avalon_jtag_slave_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_6_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_6_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave <= internal_niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave AND NOT ((niosII_system_burst_6_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_6_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave, which is an e_mux
  niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave <= (internal_niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave AND niosII_system_burst_6_downstream_read) AND NOT jtag_uart_avalon_jtag_slave_waits_for_read;
  --jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_writedata <= niosII_system_burst_6_downstream_writedata;
  --master is always granted when requested
  internal_niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave <= internal_niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave;
  --niosII_system_burst_6/downstream saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  niosII_system_burst_6_downstream_saved_grant_jtag_uart_avalon_jtag_slave <= internal_niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave;
  --allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  jtag_uart_avalon_jtag_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  jtag_uart_avalon_jtag_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  jtag_uart_avalon_jtag_slave_master_qreq_vector <= std_logic'('1');
  --jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_reset_n <= reset_n;
  jtag_uart_avalon_jtag_slave_chipselect <= internal_niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_firsttransfer <= A_WE_StdLogic((std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1'), jtag_uart_avalon_jtag_slave_unreg_firsttransfer, jtag_uart_avalon_jtag_slave_reg_firsttransfer);
  --jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_unreg_firsttransfer <= NOT ((jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND jtag_uart_avalon_jtag_slave_any_continuerequest));
  --jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1' then 
        jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  jtag_uart_avalon_jtag_slave_beginbursttransfer_internal <= jtag_uart_avalon_jtag_slave_begins_xfer;
  --~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_read_n <= NOT ((internal_niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave AND niosII_system_burst_6_downstream_read));
  --~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_write_n <= NOT ((internal_niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave AND niosII_system_burst_6_downstream_write));
  --jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_address <= niosII_system_burst_6_downstream_nativeaddress(0);
  --d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_read <= jtag_uart_avalon_jtag_slave_in_a_read_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_read_cycle <= internal_niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave AND niosII_system_burst_6_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  --jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_write <= jtag_uart_avalon_jtag_slave_in_a_write_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_write_cycle <= internal_niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave AND niosII_system_burst_6_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wait_for_jtag_uart_avalon_jtag_slave_counter <= std_logic'('0');
  --assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_irq_from_sa <= jtag_uart_avalon_jtag_slave_irq;
  --vhdl renameroo for output signals
  jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave <= internal_niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave <= internal_niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave <= internal_niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave;
--synthesis translate_off
    --jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_6/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line19 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_6_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line19, now);
          write(write_line19, string'(": "));
          write(write_line19, string'("niosII_system_burst_6/downstream drove 0 on its 'arbitrationshare' port while accessing slave jtag_uart/avalon_jtag_slave"));
          write(output, write_line19.all);
          deallocate (write_line19);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_6/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line20 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_6_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line20, now);
          write(write_line20, string'(": "));
          write(write_line20, string'("niosII_system_burst_6/downstream drove 0 on its 'burstcount' port while accessing slave jtag_uart/avalon_jtag_slave"));
          write(output, write_line20.all);
          deallocate (write_line20);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity lcd_display_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_display_control_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_7_downstream_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_7_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal niosII_system_burst_7_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_byteenable : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_7_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_lcd_display_control_slave_end_xfer : OUT STD_LOGIC;
                 signal lcd_display_control_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_display_control_slave_begintransfer : OUT STD_LOGIC;
                 signal lcd_display_control_slave_read : OUT STD_LOGIC;
                 signal lcd_display_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal lcd_display_control_slave_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal lcd_display_control_slave_write : OUT STD_LOGIC;
                 signal lcd_display_control_slave_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_7_downstream_granted_lcd_display_control_slave : OUT STD_LOGIC;
                 signal niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave : OUT STD_LOGIC;
                 signal niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave : OUT STD_LOGIC;
                 signal niosII_system_burst_7_downstream_requests_lcd_display_control_slave : OUT STD_LOGIC
              );
end entity lcd_display_control_slave_arbitrator;


architecture europa of lcd_display_control_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_lcd_display_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_lcd_display_control_slave_wait_counter_eq_0 :  STD_LOGIC;
                signal internal_niosII_system_burst_7_downstream_granted_lcd_display_control_slave :  STD_LOGIC;
                signal internal_niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave :  STD_LOGIC;
                signal internal_niosII_system_burst_7_downstream_requests_lcd_display_control_slave :  STD_LOGIC;
                signal lcd_display_control_slave_allgrants :  STD_LOGIC;
                signal lcd_display_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal lcd_display_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal lcd_display_control_slave_any_continuerequest :  STD_LOGIC;
                signal lcd_display_control_slave_arb_counter_enable :  STD_LOGIC;
                signal lcd_display_control_slave_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal lcd_display_control_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal lcd_display_control_slave_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal lcd_display_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal lcd_display_control_slave_begins_xfer :  STD_LOGIC;
                signal lcd_display_control_slave_counter_load_value :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal lcd_display_control_slave_end_xfer :  STD_LOGIC;
                signal lcd_display_control_slave_firsttransfer :  STD_LOGIC;
                signal lcd_display_control_slave_grant_vector :  STD_LOGIC;
                signal lcd_display_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal lcd_display_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal lcd_display_control_slave_master_qreq_vector :  STD_LOGIC;
                signal lcd_display_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal lcd_display_control_slave_pretend_byte_enable :  STD_LOGIC;
                signal lcd_display_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal lcd_display_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal lcd_display_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal lcd_display_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal lcd_display_control_slave_wait_counter :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal lcd_display_control_slave_waits_for_read :  STD_LOGIC;
                signal lcd_display_control_slave_waits_for_write :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_saved_grant_lcd_display_control_slave :  STD_LOGIC;
                signal wait_for_lcd_display_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT lcd_display_control_slave_end_xfer;
    end if;

  end process;

  lcd_display_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave);
  --assign lcd_display_control_slave_readdata_from_sa = lcd_display_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_display_control_slave_readdata_from_sa <= lcd_display_control_slave_readdata;
  internal_niosII_system_burst_7_downstream_requests_lcd_display_control_slave <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_7_downstream_read OR niosII_system_burst_7_downstream_write)))))));
  --lcd_display_control_slave_arb_share_counter set values, which is an e_mux
  lcd_display_control_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_7_downstream_granted_lcd_display_control_slave)) = '1'), (std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_7_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 6);
  --lcd_display_control_slave_non_bursting_master_requests mux, which is an e_mux
  lcd_display_control_slave_non_bursting_master_requests <= std_logic'('0');
  --lcd_display_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  lcd_display_control_slave_any_bursting_master_saved_grant <= niosII_system_burst_7_downstream_saved_grant_lcd_display_control_slave;
  --lcd_display_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  lcd_display_control_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(lcd_display_control_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (lcd_display_control_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(lcd_display_control_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (lcd_display_control_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --lcd_display_control_slave_allgrants all slave grants, which is an e_mux
  lcd_display_control_slave_allgrants <= lcd_display_control_slave_grant_vector;
  --lcd_display_control_slave_end_xfer assignment, which is an e_assign
  lcd_display_control_slave_end_xfer <= NOT ((lcd_display_control_slave_waits_for_read OR lcd_display_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_lcd_display_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_lcd_display_control_slave <= lcd_display_control_slave_end_xfer AND (((NOT lcd_display_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --lcd_display_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  lcd_display_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_lcd_display_control_slave AND lcd_display_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_lcd_display_control_slave AND NOT lcd_display_control_slave_non_bursting_master_requests));
  --lcd_display_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_display_control_slave_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_display_control_slave_arb_counter_enable) = '1' then 
        lcd_display_control_slave_arb_share_counter <= lcd_display_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --lcd_display_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_display_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((lcd_display_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_lcd_display_control_slave)) OR ((end_xfer_arb_share_counter_term_lcd_display_control_slave AND NOT lcd_display_control_slave_non_bursting_master_requests)))) = '1' then 
        lcd_display_control_slave_slavearbiterlockenable <= or_reduce(lcd_display_control_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_7/downstream lcd_display/control_slave arbiterlock, which is an e_assign
  niosII_system_burst_7_downstream_arbiterlock <= lcd_display_control_slave_slavearbiterlockenable AND niosII_system_burst_7_downstream_continuerequest;
  --lcd_display_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  lcd_display_control_slave_slavearbiterlockenable2 <= or_reduce(lcd_display_control_slave_arb_share_counter_next_value);
  --niosII_system_burst_7/downstream lcd_display/control_slave arbiterlock2, which is an e_assign
  niosII_system_burst_7_downstream_arbiterlock2 <= lcd_display_control_slave_slavearbiterlockenable2 AND niosII_system_burst_7_downstream_continuerequest;
  --lcd_display_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  lcd_display_control_slave_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_7_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_7_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave <= internal_niosII_system_burst_7_downstream_requests_lcd_display_control_slave AND NOT ((niosII_system_burst_7_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_7_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave, which is an e_mux
  niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave <= (internal_niosII_system_burst_7_downstream_granted_lcd_display_control_slave AND niosII_system_burst_7_downstream_read) AND NOT lcd_display_control_slave_waits_for_read;
  --lcd_display_control_slave_writedata mux, which is an e_mux
  lcd_display_control_slave_writedata <= niosII_system_burst_7_downstream_writedata;
  --master is always granted when requested
  internal_niosII_system_burst_7_downstream_granted_lcd_display_control_slave <= internal_niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave;
  --niosII_system_burst_7/downstream saved-grant lcd_display/control_slave, which is an e_assign
  niosII_system_burst_7_downstream_saved_grant_lcd_display_control_slave <= internal_niosII_system_burst_7_downstream_requests_lcd_display_control_slave;
  --allow new arb cycle for lcd_display/control_slave, which is an e_assign
  lcd_display_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  lcd_display_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  lcd_display_control_slave_master_qreq_vector <= std_logic'('1');
  lcd_display_control_slave_begintransfer <= lcd_display_control_slave_begins_xfer;
  --lcd_display_control_slave_firsttransfer first transaction, which is an e_assign
  lcd_display_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(lcd_display_control_slave_begins_xfer) = '1'), lcd_display_control_slave_unreg_firsttransfer, lcd_display_control_slave_reg_firsttransfer);
  --lcd_display_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  lcd_display_control_slave_unreg_firsttransfer <= NOT ((lcd_display_control_slave_slavearbiterlockenable AND lcd_display_control_slave_any_continuerequest));
  --lcd_display_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_display_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_display_control_slave_begins_xfer) = '1' then 
        lcd_display_control_slave_reg_firsttransfer <= lcd_display_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --lcd_display_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  lcd_display_control_slave_beginbursttransfer_internal <= lcd_display_control_slave_begins_xfer;
  --lcd_display_control_slave_read assignment, which is an e_mux
  lcd_display_control_slave_read <= (((internal_niosII_system_burst_7_downstream_granted_lcd_display_control_slave AND niosII_system_burst_7_downstream_read)) AND NOT lcd_display_control_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("0000000000000000000000000") & (lcd_display_control_slave_wait_counter))<std_logic_vector'("00000000000000000000000000011001"))));
  --lcd_display_control_slave_write assignment, which is an e_mux
  lcd_display_control_slave_write <= (((((internal_niosII_system_burst_7_downstream_granted_lcd_display_control_slave AND niosII_system_burst_7_downstream_write)) AND NOT lcd_display_control_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("0000000000000000000000000") & (lcd_display_control_slave_wait_counter))>=std_logic_vector'("00000000000000000000000000011001"))))) AND to_std_logic((((std_logic_vector'("0000000000000000000000000") & (lcd_display_control_slave_wait_counter))<std_logic_vector'("00000000000000000000000000110010"))))) AND lcd_display_control_slave_pretend_byte_enable;
  --lcd_display_control_slave_address mux, which is an e_mux
  lcd_display_control_slave_address <= niosII_system_burst_7_downstream_nativeaddress;
  --d1_lcd_display_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_lcd_display_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_lcd_display_control_slave_end_xfer <= lcd_display_control_slave_end_xfer;
    end if;

  end process;

  --lcd_display_control_slave_waits_for_read in a cycle, which is an e_mux
  lcd_display_control_slave_waits_for_read <= lcd_display_control_slave_in_a_read_cycle AND wait_for_lcd_display_control_slave_counter;
  --lcd_display_control_slave_in_a_read_cycle assignment, which is an e_assign
  lcd_display_control_slave_in_a_read_cycle <= internal_niosII_system_burst_7_downstream_granted_lcd_display_control_slave AND niosII_system_burst_7_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= lcd_display_control_slave_in_a_read_cycle;
  --lcd_display_control_slave_waits_for_write in a cycle, which is an e_mux
  lcd_display_control_slave_waits_for_write <= lcd_display_control_slave_in_a_write_cycle AND wait_for_lcd_display_control_slave_counter;
  --lcd_display_control_slave_in_a_write_cycle assignment, which is an e_assign
  lcd_display_control_slave_in_a_write_cycle <= internal_niosII_system_burst_7_downstream_granted_lcd_display_control_slave AND niosII_system_burst_7_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= lcd_display_control_slave_in_a_write_cycle;
  internal_lcd_display_control_slave_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("0000000000000000000000000") & (lcd_display_control_slave_wait_counter)) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_display_control_slave_wait_counter <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      lcd_display_control_slave_wait_counter <= lcd_display_control_slave_counter_load_value;
    end if;

  end process;

  lcd_display_control_slave_counter_load_value <= A_EXT (A_WE_StdLogicVector((std_logic'(((lcd_display_control_slave_in_a_write_cycle AND lcd_display_control_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000001001001"), A_WE_StdLogicVector((std_logic'(((lcd_display_control_slave_in_a_read_cycle AND lcd_display_control_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000110000"), A_WE_StdLogicVector((std_logic'((NOT internal_lcd_display_control_slave_wait_counter_eq_0)) = '1'), ((std_logic_vector'("00000000000000000000000000") & (lcd_display_control_slave_wait_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000")))), 7);
  wait_for_lcd_display_control_slave_counter <= lcd_display_control_slave_begins_xfer OR NOT internal_lcd_display_control_slave_wait_counter_eq_0;
  --lcd_display_control_slave_pretend_byte_enable byte enable port mux, which is an e_mux
  lcd_display_control_slave_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_7_downstream_granted_lcd_display_control_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_7_downstream_byteenable))), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  lcd_display_control_slave_wait_counter_eq_0 <= internal_lcd_display_control_slave_wait_counter_eq_0;
  --vhdl renameroo for output signals
  niosII_system_burst_7_downstream_granted_lcd_display_control_slave <= internal_niosII_system_burst_7_downstream_granted_lcd_display_control_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave <= internal_niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_7_downstream_requests_lcd_display_control_slave <= internal_niosII_system_burst_7_downstream_requests_lcd_display_control_slave;
--synthesis translate_off
    --lcd_display/control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_7/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line21 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_7_downstream_requests_lcd_display_control_slave AND to_std_logic((((std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_7_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line21, now);
          write(write_line21, string'(": "));
          write(write_line21, string'("niosII_system_burst_7/downstream drove 0 on its 'arbitrationshare' port while accessing slave lcd_display/control_slave"));
          write(output, write_line21.all);
          deallocate (write_line21);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_7/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line22 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_7_downstream_requests_lcd_display_control_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_7_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line22, now);
          write(write_line22, string'(": "));
          write(write_line22, string'("niosII_system_burst_7/downstream drove 0 on its 'burstcount' port while accessing slave lcd_display/control_slave"));
          write(output, write_line22.all);
          deallocate (write_line22);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity led_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal led_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_8_downstream_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_8_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal niosII_system_burst_8_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_byteenable : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_8_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_led_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal led_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal led_pio_s1_chipselect : OUT STD_LOGIC;
                 signal led_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal led_pio_s1_reset_n : OUT STD_LOGIC;
                 signal led_pio_s1_write_n : OUT STD_LOGIC;
                 signal led_pio_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_8_downstream_granted_led_pio_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_8_downstream_qualified_request_led_pio_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_8_downstream_read_data_valid_led_pio_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_8_downstream_requests_led_pio_s1 : OUT STD_LOGIC
              );
end entity led_pio_s1_arbitrator;


architecture europa of led_pio_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_led_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_8_downstream_granted_led_pio_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_8_downstream_qualified_request_led_pio_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_8_downstream_requests_led_pio_s1 :  STD_LOGIC;
                signal led_pio_s1_allgrants :  STD_LOGIC;
                signal led_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal led_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal led_pio_s1_any_continuerequest :  STD_LOGIC;
                signal led_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal led_pio_s1_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal led_pio_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal led_pio_s1_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal led_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal led_pio_s1_begins_xfer :  STD_LOGIC;
                signal led_pio_s1_end_xfer :  STD_LOGIC;
                signal led_pio_s1_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_grant_vector :  STD_LOGIC;
                signal led_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal led_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal led_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal led_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal led_pio_s1_pretend_byte_enable :  STD_LOGIC;
                signal led_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal led_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal led_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_waits_for_read :  STD_LOGIC;
                signal led_pio_s1_waits_for_write :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_saved_grant_led_pio_s1 :  STD_LOGIC;
                signal wait_for_led_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT led_pio_s1_end_xfer;
    end if;

  end process;

  led_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_8_downstream_qualified_request_led_pio_s1);
  --assign led_pio_s1_readdata_from_sa = led_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  led_pio_s1_readdata_from_sa <= led_pio_s1_readdata;
  internal_niosII_system_burst_8_downstream_requests_led_pio_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_8_downstream_read OR niosII_system_burst_8_downstream_write)))))));
  --led_pio_s1_arb_share_counter set values, which is an e_mux
  led_pio_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_8_downstream_granted_led_pio_s1)) = '1'), (std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_8_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 6);
  --led_pio_s1_non_bursting_master_requests mux, which is an e_mux
  led_pio_s1_non_bursting_master_requests <= std_logic'('0');
  --led_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  led_pio_s1_any_bursting_master_saved_grant <= niosII_system_burst_8_downstream_saved_grant_led_pio_s1;
  --led_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  led_pio_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(led_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (led_pio_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(led_pio_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (led_pio_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --led_pio_s1_allgrants all slave grants, which is an e_mux
  led_pio_s1_allgrants <= led_pio_s1_grant_vector;
  --led_pio_s1_end_xfer assignment, which is an e_assign
  led_pio_s1_end_xfer <= NOT ((led_pio_s1_waits_for_read OR led_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_led_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_led_pio_s1 <= led_pio_s1_end_xfer AND (((NOT led_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --led_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  led_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_led_pio_s1 AND led_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_led_pio_s1 AND NOT led_pio_s1_non_bursting_master_requests));
  --led_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(led_pio_s1_arb_counter_enable) = '1' then 
        led_pio_s1_arb_share_counter <= led_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --led_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((led_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_led_pio_s1)) OR ((end_xfer_arb_share_counter_term_led_pio_s1 AND NOT led_pio_s1_non_bursting_master_requests)))) = '1' then 
        led_pio_s1_slavearbiterlockenable <= or_reduce(led_pio_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_8/downstream led_pio/s1 arbiterlock, which is an e_assign
  niosII_system_burst_8_downstream_arbiterlock <= led_pio_s1_slavearbiterlockenable AND niosII_system_burst_8_downstream_continuerequest;
  --led_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  led_pio_s1_slavearbiterlockenable2 <= or_reduce(led_pio_s1_arb_share_counter_next_value);
  --niosII_system_burst_8/downstream led_pio/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_8_downstream_arbiterlock2 <= led_pio_s1_slavearbiterlockenable2 AND niosII_system_burst_8_downstream_continuerequest;
  --led_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  led_pio_s1_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_8_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_8_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_8_downstream_qualified_request_led_pio_s1 <= internal_niosII_system_burst_8_downstream_requests_led_pio_s1 AND NOT ((niosII_system_burst_8_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_8_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_8_downstream_read_data_valid_led_pio_s1, which is an e_mux
  niosII_system_burst_8_downstream_read_data_valid_led_pio_s1 <= (internal_niosII_system_burst_8_downstream_granted_led_pio_s1 AND niosII_system_burst_8_downstream_read) AND NOT led_pio_s1_waits_for_read;
  --led_pio_s1_writedata mux, which is an e_mux
  led_pio_s1_writedata <= niosII_system_burst_8_downstream_writedata;
  --master is always granted when requested
  internal_niosII_system_burst_8_downstream_granted_led_pio_s1 <= internal_niosII_system_burst_8_downstream_qualified_request_led_pio_s1;
  --niosII_system_burst_8/downstream saved-grant led_pio/s1, which is an e_assign
  niosII_system_burst_8_downstream_saved_grant_led_pio_s1 <= internal_niosII_system_burst_8_downstream_requests_led_pio_s1;
  --allow new arb cycle for led_pio/s1, which is an e_assign
  led_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  led_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  led_pio_s1_master_qreq_vector <= std_logic'('1');
  --led_pio_s1_reset_n assignment, which is an e_assign
  led_pio_s1_reset_n <= reset_n;
  led_pio_s1_chipselect <= internal_niosII_system_burst_8_downstream_granted_led_pio_s1;
  --led_pio_s1_firsttransfer first transaction, which is an e_assign
  led_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(led_pio_s1_begins_xfer) = '1'), led_pio_s1_unreg_firsttransfer, led_pio_s1_reg_firsttransfer);
  --led_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  led_pio_s1_unreg_firsttransfer <= NOT ((led_pio_s1_slavearbiterlockenable AND led_pio_s1_any_continuerequest));
  --led_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(led_pio_s1_begins_xfer) = '1' then 
        led_pio_s1_reg_firsttransfer <= led_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --led_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  led_pio_s1_beginbursttransfer_internal <= led_pio_s1_begins_xfer;
  --~led_pio_s1_write_n assignment, which is an e_mux
  led_pio_s1_write_n <= NOT ((((internal_niosII_system_burst_8_downstream_granted_led_pio_s1 AND niosII_system_burst_8_downstream_write)) AND led_pio_s1_pretend_byte_enable));
  --led_pio_s1_address mux, which is an e_mux
  led_pio_s1_address <= niosII_system_burst_8_downstream_nativeaddress;
  --d1_led_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_led_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_led_pio_s1_end_xfer <= led_pio_s1_end_xfer;
    end if;

  end process;

  --led_pio_s1_waits_for_read in a cycle, which is an e_mux
  led_pio_s1_waits_for_read <= led_pio_s1_in_a_read_cycle AND led_pio_s1_begins_xfer;
  --led_pio_s1_in_a_read_cycle assignment, which is an e_assign
  led_pio_s1_in_a_read_cycle <= internal_niosII_system_burst_8_downstream_granted_led_pio_s1 AND niosII_system_burst_8_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= led_pio_s1_in_a_read_cycle;
  --led_pio_s1_waits_for_write in a cycle, which is an e_mux
  led_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --led_pio_s1_in_a_write_cycle assignment, which is an e_assign
  led_pio_s1_in_a_write_cycle <= internal_niosII_system_burst_8_downstream_granted_led_pio_s1 AND niosII_system_burst_8_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= led_pio_s1_in_a_write_cycle;
  wait_for_led_pio_s1_counter <= std_logic'('0');
  --led_pio_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  led_pio_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_8_downstream_granted_led_pio_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_8_downstream_byteenable))), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  niosII_system_burst_8_downstream_granted_led_pio_s1 <= internal_niosII_system_burst_8_downstream_granted_led_pio_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_8_downstream_qualified_request_led_pio_s1 <= internal_niosII_system_burst_8_downstream_qualified_request_led_pio_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_8_downstream_requests_led_pio_s1 <= internal_niosII_system_burst_8_downstream_requests_led_pio_s1;
--synthesis translate_off
    --led_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_8/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line23 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_8_downstream_requests_led_pio_s1 AND to_std_logic((((std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_8_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line23, now);
          write(write_line23, string'(": "));
          write(write_line23, string'("niosII_system_burst_8/downstream drove 0 on its 'arbitrationshare' port while accessing slave led_pio/s1"));
          write(output, write_line23.all);
          deallocate (write_line23);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_8/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line24 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_8_downstream_requests_led_pio_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_8_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line24, now);
          write(write_line24, string'(": "));
          write(write_line24, string'("niosII_system_burst_8/downstream drove 0 on its 'burstcount' port while accessing slave led_pio/s1"));
          write(output, write_line24.all);
          deallocate (write_line24);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity memory_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_2_downstream_address_to_slave : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal niosII_system_burst_2_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_2_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_2_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_3_downstream_address_to_slave : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal niosII_system_burst_3_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_3_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_3_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_memory_s1_end_xfer : OUT STD_LOGIC;
                 signal memory_s1_address : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal memory_s1_chipselect : OUT STD_LOGIC;
                 signal memory_s1_clken : OUT STD_LOGIC;
                 signal memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal memory_s1_reset : OUT STD_LOGIC;
                 signal memory_s1_write : OUT STD_LOGIC;
                 signal memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_2_downstream_granted_memory_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_2_downstream_qualified_request_memory_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_2_downstream_read_data_valid_memory_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_2_downstream_requests_memory_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_3_downstream_granted_memory_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_3_downstream_qualified_request_memory_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_3_downstream_read_data_valid_memory_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_3_downstream_requests_memory_s1 : OUT STD_LOGIC
              );
end entity memory_s1_arbitrator;


architecture europa of memory_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_memory_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_2_downstream_granted_memory_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_2_downstream_qualified_request_memory_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_2_downstream_requests_memory_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_3_downstream_granted_memory_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_3_downstream_qualified_request_memory_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_3_downstream_requests_memory_s1 :  STD_LOGIC;
                signal last_cycle_niosII_system_burst_2_downstream_granted_slave_memory_s1 :  STD_LOGIC;
                signal last_cycle_niosII_system_burst_3_downstream_granted_slave_memory_s1 :  STD_LOGIC;
                signal memory_s1_allgrants :  STD_LOGIC;
                signal memory_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal memory_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal memory_s1_any_continuerequest :  STD_LOGIC;
                signal memory_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal memory_s1_arb_counter_enable :  STD_LOGIC;
                signal memory_s1_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal memory_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal memory_s1_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal memory_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal memory_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal memory_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal memory_s1_begins_xfer :  STD_LOGIC;
                signal memory_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal memory_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal memory_s1_end_xfer :  STD_LOGIC;
                signal memory_s1_firsttransfer :  STD_LOGIC;
                signal memory_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal memory_s1_in_a_read_cycle :  STD_LOGIC;
                signal memory_s1_in_a_write_cycle :  STD_LOGIC;
                signal memory_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal memory_s1_non_bursting_master_requests :  STD_LOGIC;
                signal memory_s1_reg_firsttransfer :  STD_LOGIC;
                signal memory_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal memory_s1_slavearbiterlockenable :  STD_LOGIC;
                signal memory_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal memory_s1_unreg_firsttransfer :  STD_LOGIC;
                signal memory_s1_waits_for_read :  STD_LOGIC;
                signal memory_s1_waits_for_write :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register_in :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_saved_grant_memory_s1 :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register_in :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_saved_grant_memory_s1 :  STD_LOGIC;
                signal p1_niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register :  STD_LOGIC;
                signal p1_niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register :  STD_LOGIC;
                signal shifted_address_to_memory_s1_from_niosII_system_burst_2_downstream :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal shifted_address_to_memory_s1_from_niosII_system_burst_3_downstream :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal wait_for_memory_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT memory_s1_end_xfer;
    end if;

  end process;

  memory_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_niosII_system_burst_2_downstream_qualified_request_memory_s1 OR internal_niosII_system_burst_3_downstream_qualified_request_memory_s1));
  --assign memory_s1_readdata_from_sa = memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  memory_s1_readdata_from_sa <= memory_s1_readdata;
  internal_niosII_system_burst_2_downstream_requests_memory_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_2_downstream_read OR niosII_system_burst_2_downstream_write)))))));
  --memory_s1_arb_share_counter set values, which is an e_mux
  memory_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_2_downstream_granted_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_2_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_3_downstream_granted_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_3_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_2_downstream_granted_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_2_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_3_downstream_granted_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_3_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001"))))), 4);
  --memory_s1_non_bursting_master_requests mux, which is an e_mux
  memory_s1_non_bursting_master_requests <= std_logic'('0');
  --memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  memory_s1_any_bursting_master_saved_grant <= ((niosII_system_burst_2_downstream_saved_grant_memory_s1 OR niosII_system_burst_3_downstream_saved_grant_memory_s1) OR niosII_system_burst_2_downstream_saved_grant_memory_s1) OR niosII_system_burst_3_downstream_saved_grant_memory_s1;
  --memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  memory_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(memory_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (memory_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(memory_s1_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (memory_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --memory_s1_allgrants all slave grants, which is an e_mux
  memory_s1_allgrants <= (((or_reduce(memory_s1_grant_vector)) OR (or_reduce(memory_s1_grant_vector))) OR (or_reduce(memory_s1_grant_vector))) OR (or_reduce(memory_s1_grant_vector));
  --memory_s1_end_xfer assignment, which is an e_assign
  memory_s1_end_xfer <= NOT ((memory_s1_waits_for_read OR memory_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_memory_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_memory_s1 <= memory_s1_end_xfer AND (((NOT memory_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  memory_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_memory_s1 AND memory_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_memory_s1 AND NOT memory_s1_non_bursting_master_requests));
  --memory_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      memory_s1_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(memory_s1_arb_counter_enable) = '1' then 
        memory_s1_arb_share_counter <= memory_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      memory_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(memory_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_memory_s1)) OR ((end_xfer_arb_share_counter_term_memory_s1 AND NOT memory_s1_non_bursting_master_requests)))) = '1' then 
        memory_s1_slavearbiterlockenable <= or_reduce(memory_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_2/downstream memory/s1 arbiterlock, which is an e_assign
  niosII_system_burst_2_downstream_arbiterlock <= memory_s1_slavearbiterlockenable AND niosII_system_burst_2_downstream_continuerequest;
  --memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  memory_s1_slavearbiterlockenable2 <= or_reduce(memory_s1_arb_share_counter_next_value);
  --niosII_system_burst_2/downstream memory/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_2_downstream_arbiterlock2 <= memory_s1_slavearbiterlockenable2 AND niosII_system_burst_2_downstream_continuerequest;
  --niosII_system_burst_3/downstream memory/s1 arbiterlock, which is an e_assign
  niosII_system_burst_3_downstream_arbiterlock <= memory_s1_slavearbiterlockenable AND niosII_system_burst_3_downstream_continuerequest;
  --niosII_system_burst_3/downstream memory/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_3_downstream_arbiterlock2 <= memory_s1_slavearbiterlockenable2 AND niosII_system_burst_3_downstream_continuerequest;
  --niosII_system_burst_3/downstream granted memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_niosII_system_burst_3_downstream_granted_slave_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_niosII_system_burst_3_downstream_granted_slave_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(niosII_system_burst_3_downstream_saved_grant_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(memory_s1_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_3_downstream_granted_slave_memory_s1))))));
    end if;

  end process;

  --niosII_system_burst_3_downstream_continuerequest continued request, which is an e_mux
  niosII_system_burst_3_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_3_downstream_granted_slave_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --memory_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  memory_s1_any_continuerequest <= niosII_system_burst_3_downstream_continuerequest OR niosII_system_burst_2_downstream_continuerequest;
  internal_niosII_system_burst_2_downstream_qualified_request_memory_s1 <= internal_niosII_system_burst_2_downstream_requests_memory_s1 AND NOT (niosII_system_burst_3_downstream_arbiterlock);
  --niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register_in <= (internal_niosII_system_burst_2_downstream_granted_memory_s1 AND niosII_system_burst_2_downstream_read) AND NOT memory_s1_waits_for_read;
  --shift register p1 niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register) & A_ToStdLogicVector(niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register_in)));
  --niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register <= p1_niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid niosII_system_burst_2_downstream_read_data_valid_memory_s1, which is an e_mux
  niosII_system_burst_2_downstream_read_data_valid_memory_s1 <= niosII_system_burst_2_downstream_read_data_valid_memory_s1_shift_register;
  --memory_s1_writedata mux, which is an e_mux
  memory_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_2_downstream_granted_memory_s1)) = '1'), niosII_system_burst_2_downstream_writedata, niosII_system_burst_3_downstream_writedata);
  --mux memory_s1_clken, which is an e_mux
  memory_s1_clken <= std_logic'('1');
  internal_niosII_system_burst_3_downstream_requests_memory_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_3_downstream_read OR niosII_system_burst_3_downstream_write)))))));
  --niosII_system_burst_2/downstream granted memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_niosII_system_burst_2_downstream_granted_slave_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_niosII_system_burst_2_downstream_granted_slave_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(niosII_system_burst_2_downstream_saved_grant_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(memory_s1_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_2_downstream_granted_slave_memory_s1))))));
    end if;

  end process;

  --niosII_system_burst_2_downstream_continuerequest continued request, which is an e_mux
  niosII_system_burst_2_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_2_downstream_granted_slave_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  internal_niosII_system_burst_3_downstream_qualified_request_memory_s1 <= internal_niosII_system_burst_3_downstream_requests_memory_s1 AND NOT (niosII_system_burst_2_downstream_arbiterlock);
  --niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register_in <= (internal_niosII_system_burst_3_downstream_granted_memory_s1 AND niosII_system_burst_3_downstream_read) AND NOT memory_s1_waits_for_read;
  --shift register p1 niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register) & A_ToStdLogicVector(niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register_in)));
  --niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register <= p1_niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid niosII_system_burst_3_downstream_read_data_valid_memory_s1, which is an e_mux
  niosII_system_burst_3_downstream_read_data_valid_memory_s1 <= niosII_system_burst_3_downstream_read_data_valid_memory_s1_shift_register;
  --allow new arb cycle for memory/s1, which is an e_assign
  memory_s1_allow_new_arb_cycle <= NOT niosII_system_burst_2_downstream_arbiterlock AND NOT niosII_system_burst_3_downstream_arbiterlock;
  --niosII_system_burst_3/downstream assignment into master qualified-requests vector for memory/s1, which is an e_assign
  memory_s1_master_qreq_vector(0) <= internal_niosII_system_burst_3_downstream_qualified_request_memory_s1;
  --niosII_system_burst_3/downstream grant memory/s1, which is an e_assign
  internal_niosII_system_burst_3_downstream_granted_memory_s1 <= memory_s1_grant_vector(0);
  --niosII_system_burst_3/downstream saved-grant memory/s1, which is an e_assign
  niosII_system_burst_3_downstream_saved_grant_memory_s1 <= memory_s1_arb_winner(0);
  --niosII_system_burst_2/downstream assignment into master qualified-requests vector for memory/s1, which is an e_assign
  memory_s1_master_qreq_vector(1) <= internal_niosII_system_burst_2_downstream_qualified_request_memory_s1;
  --niosII_system_burst_2/downstream grant memory/s1, which is an e_assign
  internal_niosII_system_burst_2_downstream_granted_memory_s1 <= memory_s1_grant_vector(1);
  --niosII_system_burst_2/downstream saved-grant memory/s1, which is an e_assign
  niosII_system_burst_2_downstream_saved_grant_memory_s1 <= memory_s1_arb_winner(1);
  --memory/s1 chosen-master double-vector, which is an e_assign
  memory_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((memory_s1_master_qreq_vector & memory_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT memory_s1_master_qreq_vector & NOT memory_s1_master_qreq_vector))) + (std_logic_vector'("000") & (memory_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  memory_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((memory_s1_allow_new_arb_cycle AND or_reduce(memory_s1_grant_vector)))) = '1'), memory_s1_grant_vector, memory_s1_saved_chosen_master_vector);
  --saved memory_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      memory_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(memory_s1_allow_new_arb_cycle) = '1' then 
        memory_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(memory_s1_grant_vector)) = '1'), memory_s1_grant_vector, memory_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  memory_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((memory_s1_chosen_master_double_vector(1) OR memory_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((memory_s1_chosen_master_double_vector(0) OR memory_s1_chosen_master_double_vector(2)))));
  --memory/s1 chosen master rotated left, which is an e_assign
  memory_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(memory_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(memory_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --memory/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      memory_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(memory_s1_grant_vector)) = '1' then 
        memory_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(memory_s1_end_xfer) = '1'), memory_s1_chosen_master_rot_left, memory_s1_grant_vector);
      end if;
    end if;

  end process;

  --~memory_s1_reset assignment, which is an e_assign
  memory_s1_reset <= NOT reset_n;
  memory_s1_chipselect <= internal_niosII_system_burst_2_downstream_granted_memory_s1 OR internal_niosII_system_burst_3_downstream_granted_memory_s1;
  --memory_s1_firsttransfer first transaction, which is an e_assign
  memory_s1_firsttransfer <= A_WE_StdLogic((std_logic'(memory_s1_begins_xfer) = '1'), memory_s1_unreg_firsttransfer, memory_s1_reg_firsttransfer);
  --memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  memory_s1_unreg_firsttransfer <= NOT ((memory_s1_slavearbiterlockenable AND memory_s1_any_continuerequest));
  --memory_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      memory_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(memory_s1_begins_xfer) = '1' then 
        memory_s1_reg_firsttransfer <= memory_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  memory_s1_beginbursttransfer_internal <= memory_s1_begins_xfer;
  --memory_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  memory_s1_arbitration_holdoff_internal <= memory_s1_begins_xfer AND memory_s1_firsttransfer;
  --memory_s1_write assignment, which is an e_mux
  memory_s1_write <= ((internal_niosII_system_burst_2_downstream_granted_memory_s1 AND niosII_system_burst_2_downstream_write)) OR ((internal_niosII_system_burst_3_downstream_granted_memory_s1 AND niosII_system_burst_3_downstream_write));
  shifted_address_to_memory_s1_from_niosII_system_burst_2_downstream <= niosII_system_burst_2_downstream_address_to_slave;
  --memory_s1_address mux, which is an e_mux
  memory_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_2_downstream_granted_memory_s1)) = '1'), (A_SRL(shifted_address_to_memory_s1_from_niosII_system_burst_2_downstream,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_memory_s1_from_niosII_system_burst_3_downstream,std_logic_vector'("00000000000000000000000000000010")))), 12);
  shifted_address_to_memory_s1_from_niosII_system_burst_3_downstream <= niosII_system_burst_3_downstream_address_to_slave;
  --d1_memory_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_memory_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_memory_s1_end_xfer <= memory_s1_end_xfer;
    end if;

  end process;

  --memory_s1_waits_for_read in a cycle, which is an e_mux
  memory_s1_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(memory_s1_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --memory_s1_in_a_read_cycle assignment, which is an e_assign
  memory_s1_in_a_read_cycle <= ((internal_niosII_system_burst_2_downstream_granted_memory_s1 AND niosII_system_burst_2_downstream_read)) OR ((internal_niosII_system_burst_3_downstream_granted_memory_s1 AND niosII_system_burst_3_downstream_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= memory_s1_in_a_read_cycle;
  --memory_s1_waits_for_write in a cycle, which is an e_mux
  memory_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(memory_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --memory_s1_in_a_write_cycle assignment, which is an e_assign
  memory_s1_in_a_write_cycle <= ((internal_niosII_system_burst_2_downstream_granted_memory_s1 AND niosII_system_burst_2_downstream_write)) OR ((internal_niosII_system_burst_3_downstream_granted_memory_s1 AND niosII_system_burst_3_downstream_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= memory_s1_in_a_write_cycle;
  wait_for_memory_s1_counter <= std_logic'('0');
  --memory_s1_byteenable byte enable port mux, which is an e_mux
  memory_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_2_downstream_granted_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_2_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_3_downstream_granted_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_3_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  --vhdl renameroo for output signals
  niosII_system_burst_2_downstream_granted_memory_s1 <= internal_niosII_system_burst_2_downstream_granted_memory_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_2_downstream_qualified_request_memory_s1 <= internal_niosII_system_burst_2_downstream_qualified_request_memory_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_2_downstream_requests_memory_s1 <= internal_niosII_system_burst_2_downstream_requests_memory_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_3_downstream_granted_memory_s1 <= internal_niosII_system_burst_3_downstream_granted_memory_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_3_downstream_qualified_request_memory_s1 <= internal_niosII_system_burst_3_downstream_qualified_request_memory_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_3_downstream_requests_memory_s1 <= internal_niosII_system_burst_3_downstream_requests_memory_s1;
--synthesis translate_off
    --memory/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_2/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line25 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_2_downstream_requests_memory_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_2_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line25, now);
          write(write_line25, string'(": "));
          write(write_line25, string'("niosII_system_burst_2/downstream drove 0 on its 'arbitrationshare' port while accessing slave memory/s1"));
          write(output, write_line25.all);
          deallocate (write_line25);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_2/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line26 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_2_downstream_requests_memory_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_2_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line26, now);
          write(write_line26, string'(": "));
          write(write_line26, string'("niosII_system_burst_2/downstream drove 0 on its 'burstcount' port while accessing slave memory/s1"));
          write(output, write_line26.all);
          deallocate (write_line26);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_3/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line27 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_3_downstream_requests_memory_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_3_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line27, now);
          write(write_line27, string'(": "));
          write(write_line27, string'("niosII_system_burst_3/downstream drove 0 on its 'arbitrationshare' port while accessing slave memory/s1"));
          write(output, write_line27.all);
          deallocate (write_line27);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_3/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line28 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_3_downstream_requests_memory_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_3_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line28, now);
          write(write_line28, string'(": "));
          write(write_line28, string'("niosII_system_burst_3/downstream drove 0 on its 'burstcount' port while accessing slave memory/s1"));
          write(output, write_line28.all);
          deallocate (write_line28);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line29 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_2_downstream_granted_memory_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_3_downstream_granted_memory_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line29, now);
          write(write_line29, string'(": "));
          write(write_line29, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line29.all);
          deallocate (write_line29);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line30 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(niosII_system_burst_2_downstream_saved_grant_memory_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(niosII_system_burst_3_downstream_saved_grant_memory_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line30, now);
          write(write_line30, string'(": "));
          write(write_line30, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line30.all);
          deallocate (write_line30);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_0_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_0_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_0_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_0_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_0_upstream_module;


architecture europa of rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_0_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_0_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : IN STD_LOGIC;
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : IN STD_LOGIC;
                 signal niosII_system_burst_0_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_0_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_0_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_instruction_master_granted_niosII_system_burst_0_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_instruction_master_requests_niosII_system_burst_0_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_0_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_0_upstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal niosII_system_burst_0_upstream_byteaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal niosII_system_burst_0_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_0_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_0_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_0_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_0_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_0_upstream_write : OUT STD_LOGIC
              );
end entity niosII_system_burst_0_upstream_arbitrator;


architecture europa of niosII_system_burst_0_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_0_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_0_upstream_module;

component rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_0_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_0_upstream_module;

                signal cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_output_from_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal cpu_instruction_master_saved_grant_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_instruction_master_granted_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal internal_cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal internal_cpu_instruction_master_requests_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_0_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal module_input :  STD_LOGIC;
                signal module_input1 :  STD_LOGIC;
                signal module_input2 :  STD_LOGIC;
                signal module_input3 :  STD_LOGIC;
                signal module_input4 :  STD_LOGIC;
                signal module_input5 :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_0_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_0_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_0_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_0_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_0_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_0_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_0_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_0_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_0_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_0_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_0_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_0_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream);
  --assign niosII_system_burst_0_upstream_readdata_from_sa = niosII_system_burst_0_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_0_upstream_readdata_from_sa <= niosII_system_burst_0_upstream_readdata;
  internal_cpu_instruction_master_requests_niosII_system_burst_0_upstream <= ((to_std_logic(((Std_Logic_Vector'(cpu_instruction_master_address_to_slave(24 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("1100100001000100000000000")))) AND (cpu_instruction_master_read))) AND cpu_instruction_master_read;
  --assign niosII_system_burst_0_upstream_waitrequest_from_sa = niosII_system_burst_0_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_0_upstream_waitrequest_from_sa <= niosII_system_burst_0_upstream_waitrequest;
  --assign niosII_system_burst_0_upstream_readdatavalid_from_sa = niosII_system_burst_0_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_0_upstream_readdatavalid_from_sa <= niosII_system_burst_0_upstream_readdatavalid;
  --niosII_system_burst_0_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_0_upstream_arb_share_set_values <= std_logic_vector'("00000001");
  --niosII_system_burst_0_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_0_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_0_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_0_upstream_any_bursting_master_saved_grant <= cpu_instruction_master_saved_grant_niosII_system_burst_0_upstream;
  --niosII_system_burst_0_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_0_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_0_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_0_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_0_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_0_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_0_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_0_upstream_allgrants <= niosII_system_burst_0_upstream_grant_vector;
  --niosII_system_burst_0_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_0_upstream_end_xfer <= NOT ((niosII_system_burst_0_upstream_waits_for_read OR niosII_system_burst_0_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_0_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_0_upstream <= niosII_system_burst_0_upstream_end_xfer AND (((NOT niosII_system_burst_0_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_0_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_0_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_0_upstream AND niosII_system_burst_0_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_0_upstream AND NOT niosII_system_burst_0_upstream_non_bursting_master_requests));
  --niosII_system_burst_0_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_0_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_0_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_0_upstream_arb_share_counter <= niosII_system_burst_0_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_0_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_0_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_0_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_0_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_0_upstream AND NOT niosII_system_burst_0_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_0_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_0_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/instruction_master niosII_system_burst_0/upstream arbiterlock, which is an e_assign
  cpu_instruction_master_arbiterlock <= niosII_system_burst_0_upstream_slavearbiterlockenable AND cpu_instruction_master_continuerequest;
  --niosII_system_burst_0_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_0_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_0_upstream_arb_share_counter_next_value);
  --cpu/instruction_master niosII_system_burst_0/upstream arbiterlock2, which is an e_assign
  cpu_instruction_master_arbiterlock2 <= niosII_system_burst_0_upstream_slavearbiterlockenable2 AND cpu_instruction_master_continuerequest;
  --niosII_system_burst_0_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_0_upstream_any_continuerequest <= std_logic'('1');
  --cpu_instruction_master_continuerequest continued request, which is an e_assign
  cpu_instruction_master_continuerequest <= std_logic'('1');
  internal_cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_0_upstream AND NOT ((cpu_instruction_master_read AND (((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_latency_counter))))))) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register)))));
  --unique name for niosII_system_burst_0_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_0_upstream_move_on_to_next_transaction <= niosII_system_burst_0_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_0_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_0_upstream, which is an e_mux
  niosII_system_burst_0_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_niosII_system_burst_0_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_instruction_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_0_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_0_upstream : burstcount_fifo_for_niosII_system_burst_0_upstream_module
    port map(
      data_out => niosII_system_burst_0_upstream_transaction_burst_count,
      empty => niosII_system_burst_0_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input,
      clk => clk,
      data_in => niosII_system_burst_0_upstream_selected_burstcount,
      read => niosII_system_burst_0_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input1,
      write => module_input2
    );

  module_input <= std_logic'('0');
  module_input1 <= std_logic'('0');
  module_input2 <= ((in_a_read_cycle AND NOT niosII_system_burst_0_upstream_waits_for_read) AND niosII_system_burst_0_upstream_load_fifo) AND NOT ((niosII_system_burst_0_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_0_upstream_burstcount_fifo_empty));

  --niosII_system_burst_0_upstream current burst minus one, which is an e_assign
  niosII_system_burst_0_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_0_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_0_upstream, which is an e_mux
  niosII_system_burst_0_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_0_upstream_waits_for_read)) AND NOT niosII_system_burst_0_upstream_load_fifo))) = '1'), niosII_system_burst_0_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_0_upstream_waits_for_read) AND niosII_system_burst_0_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_0_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_0_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_0_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_0_upstream_transaction_burst_count, niosII_system_burst_0_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_0_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_0_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_0_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_0_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_0_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_0_upstream_current_burst <= niosII_system_burst_0_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_0_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_0_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_0_upstream_waits_for_read)) AND niosII_system_burst_0_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_0_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_0_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_0_upstream_waits_for_read)) AND NOT niosII_system_burst_0_upstream_load_fifo) OR niosII_system_burst_0_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_0_upstream_load_fifo <= p0_niosII_system_burst_0_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_0_upstream, which is an e_assign
  niosII_system_burst_0_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_0_upstream_current_burst_minus_one)) AND niosII_system_burst_0_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_0_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_0_upstream : rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_0_upstream_module
    port map(
      data_out => cpu_instruction_master_rdv_fifo_output_from_niosII_system_burst_0_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_0_upstream,
      full => open,
      clear_fifo => module_input3,
      clk => clk,
      data_in => internal_cpu_instruction_master_granted_niosII_system_burst_0_upstream,
      read => niosII_system_burst_0_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input4,
      write => module_input5
    );

  module_input3 <= std_logic'('0');
  module_input4 <= std_logic'('0');
  module_input5 <= in_a_read_cycle AND NOT niosII_system_burst_0_upstream_waits_for_read;

  cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register <= NOT cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_0_upstream;
  --local readdatavalid cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream, which is an e_mux
  cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream <= niosII_system_burst_0_upstream_readdatavalid_from_sa;
  --byteaddress mux for niosII_system_burst_0/upstream, which is an e_mux
  niosII_system_burst_0_upstream_byteaddress <= cpu_instruction_master_address_to_slave (12 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_instruction_master_granted_niosII_system_burst_0_upstream <= internal_cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream;
  --cpu/instruction_master saved-grant niosII_system_burst_0/upstream, which is an e_assign
  cpu_instruction_master_saved_grant_niosII_system_burst_0_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_0_upstream;
  --allow new arb cycle for niosII_system_burst_0/upstream, which is an e_assign
  niosII_system_burst_0_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_0_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_0_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_0_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_0_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_0_upstream_begins_xfer) = '1'), niosII_system_burst_0_upstream_unreg_firsttransfer, niosII_system_burst_0_upstream_reg_firsttransfer);
  --niosII_system_burst_0_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_0_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_0_upstream_slavearbiterlockenable AND niosII_system_burst_0_upstream_any_continuerequest));
  --niosII_system_burst_0_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_0_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_0_upstream_begins_xfer) = '1' then 
        niosII_system_burst_0_upstream_reg_firsttransfer <= niosII_system_burst_0_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_0_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_0_upstream_beginbursttransfer_internal <= niosII_system_burst_0_upstream_begins_xfer;
  --niosII_system_burst_0_upstream_read assignment, which is an e_mux
  niosII_system_burst_0_upstream_read <= internal_cpu_instruction_master_granted_niosII_system_burst_0_upstream AND cpu_instruction_master_read;
  --niosII_system_burst_0_upstream_write assignment, which is an e_mux
  niosII_system_burst_0_upstream_write <= std_logic'('0');
  --niosII_system_burst_0_upstream_address mux, which is an e_mux
  niosII_system_burst_0_upstream_address <= cpu_instruction_master_address_to_slave (10 DOWNTO 0);
  --d1_niosII_system_burst_0_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_0_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_0_upstream_end_xfer <= niosII_system_burst_0_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_0_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_0_upstream_waits_for_read <= niosII_system_burst_0_upstream_in_a_read_cycle AND internal_niosII_system_burst_0_upstream_waitrequest_from_sa;
  --niosII_system_burst_0_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_0_upstream_in_a_read_cycle <= internal_cpu_instruction_master_granted_niosII_system_burst_0_upstream AND cpu_instruction_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_0_upstream_in_a_read_cycle;
  --niosII_system_burst_0_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_0_upstream_waits_for_write <= niosII_system_burst_0_upstream_in_a_write_cycle AND internal_niosII_system_burst_0_upstream_waitrequest_from_sa;
  --niosII_system_burst_0_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_0_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_0_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_0_upstream_counter <= std_logic'('0');
  --niosII_system_burst_0_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_0_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_0_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_instruction_master_granted_niosII_system_burst_0_upstream <= internal_cpu_instruction_master_granted_niosII_system_burst_0_upstream;
  --vhdl renameroo for output signals
  cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream <= internal_cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream;
  --vhdl renameroo for output signals
  cpu_instruction_master_requests_niosII_system_burst_0_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_0_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_0_upstream_waitrequest_from_sa <= internal_niosII_system_burst_0_upstream_waitrequest_from_sa;
--synthesis translate_off
    --niosII_system_burst_0/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/instruction_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line31 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_instruction_master_requests_niosII_system_burst_0_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_instruction_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line31, now);
          write(write_line31, string'(": "));
          write(write_line31, string'("cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_0/upstream"));
          write(output, write_line31.all);
          deallocate (write_line31);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_0_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal niosII_system_burst_0_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_0_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal niosII_system_burst_0_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_0_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_0_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_0_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_0_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_0_downstream_arbitrator;


architecture europa of niosII_system_burst_0_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_0_downstream_address_to_slave :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal internal_niosII_system_burst_0_downstream_latency_counter :  STD_LOGIC;
                signal internal_niosII_system_burst_0_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_address_last_time :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_0_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_0_downstream_is_granted_some_slave :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_niosII_system_burst_0_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_niosII_system_burst_0_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module OR NOT niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module OR NOT niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module OR NOT niosII_system_burst_0_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cpu_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_0_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module OR NOT niosII_system_burst_0_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_0_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_0_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_0_downstream_address_to_slave <= niosII_system_burst_0_downstream_address;
  --niosII_system_burst_0_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_0_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_0_downstream_read_but_no_slave_selected <= (niosII_system_burst_0_downstream_read AND niosII_system_burst_0_downstream_run) AND NOT niosII_system_burst_0_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  niosII_system_burst_0_downstream_is_granted_some_slave <= niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_0_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_0_downstream_readdatavalid <= (niosII_system_burst_0_downstream_read_but_no_slave_selected OR pre_flush_niosII_system_burst_0_downstream_readdatavalid) OR niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module;
  --niosII_system_burst_0/downstream readdata mux, which is an e_mux
  niosII_system_burst_0_downstream_readdata <= cpu_jtag_debug_module_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_0_downstream_waitrequest <= NOT niosII_system_burst_0_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_niosII_system_burst_0_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_niosII_system_burst_0_downstream_latency_counter <= p1_niosII_system_burst_0_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_niosII_system_burst_0_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((niosII_system_burst_0_downstream_run AND niosII_system_burst_0_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_0_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_0_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --niosII_system_burst_0_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_0_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_0_downstream_address_to_slave <= internal_niosII_system_burst_0_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_0_downstream_latency_counter <= internal_niosII_system_burst_0_downstream_latency_counter;
  --vhdl renameroo for output signals
  niosII_system_burst_0_downstream_waitrequest <= internal_niosII_system_burst_0_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_0_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_0_downstream_address_last_time <= std_logic_vector'("00000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_0_downstream_address_last_time <= niosII_system_burst_0_downstream_address;
      end if;

    end process;

    --niosII_system_burst_0/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_0_downstream_waitrequest AND ((niosII_system_burst_0_downstream_read OR niosII_system_burst_0_downstream_write));
      end if;

    end process;

    --niosII_system_burst_0_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line32 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_0_downstream_address /= niosII_system_burst_0_downstream_address_last_time))))) = '1' then 
          write(write_line32, now);
          write(write_line32, string'(": "));
          write(write_line32, string'("niosII_system_burst_0_downstream_address did not heed wait!!!"));
          write(output, write_line32.all);
          deallocate (write_line32);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_0_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_0_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_0_downstream_burstcount_last_time <= niosII_system_burst_0_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_0_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line33 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_0_downstream_burstcount) /= std_logic'(niosII_system_burst_0_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line33, now);
          write(write_line33, string'(": "));
          write(write_line33, string'("niosII_system_burst_0_downstream_burstcount did not heed wait!!!"));
          write(output, write_line33.all);
          deallocate (write_line33);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_0_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_0_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_0_downstream_byteenable_last_time <= niosII_system_burst_0_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_0_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line34 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_0_downstream_byteenable /= niosII_system_burst_0_downstream_byteenable_last_time))))) = '1' then 
          write(write_line34, now);
          write(write_line34, string'(": "));
          write(write_line34, string'("niosII_system_burst_0_downstream_byteenable did not heed wait!!!"));
          write(output, write_line34.all);
          deallocate (write_line34);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_0_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_0_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_0_downstream_read_last_time <= niosII_system_burst_0_downstream_read;
      end if;

    end process;

    --niosII_system_burst_0_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line35 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_0_downstream_read) /= std_logic'(niosII_system_burst_0_downstream_read_last_time)))))) = '1' then 
          write(write_line35, now);
          write(write_line35, string'(": "));
          write(write_line35, string'("niosII_system_burst_0_downstream_read did not heed wait!!!"));
          write(output, write_line35.all);
          deallocate (write_line35);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_0_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_0_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_0_downstream_write_last_time <= niosII_system_burst_0_downstream_write;
      end if;

    end process;

    --niosII_system_burst_0_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line36 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_0_downstream_write) /= std_logic'(niosII_system_burst_0_downstream_write_last_time)))))) = '1' then 
          write(write_line36, now);
          write(write_line36, string'(": "));
          write(write_line36, string'("niosII_system_burst_0_downstream_write did not heed wait!!!"));
          write(output, write_line36.all);
          deallocate (write_line36);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_0_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_0_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_0_downstream_writedata_last_time <= niosII_system_burst_0_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_0_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line37 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_0_downstream_writedata /= niosII_system_burst_0_downstream_writedata_last_time)))) AND niosII_system_burst_0_downstream_write)) = '1' then 
          write(write_line37, now);
          write(write_line37, string'(": "));
          write(write_line37, string'("niosII_system_burst_0_downstream_writedata did not heed wait!!!"));
          write(output, write_line37.all);
          deallocate (write_line37);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_1_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_1_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_1_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_1_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_1_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_1_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_1_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_1_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_1_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_1_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_1_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_1_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_1_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_1_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_1_upstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal niosII_system_burst_1_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_1_upstream_byteaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal niosII_system_burst_1_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_1_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_1_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_1_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_1_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_1_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_1_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity niosII_system_burst_1_upstream_arbitrator;


architecture europa of niosII_system_burst_1_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_1_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_1_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_1_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_1_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_1_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_1_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_1_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_1_upstream_write :  STD_LOGIC;
                signal module_input10 :  STD_LOGIC;
                signal module_input11 :  STD_LOGIC;
                signal module_input6 :  STD_LOGIC;
                signal module_input7 :  STD_LOGIC;
                signal module_input8 :  STD_LOGIC;
                signal module_input9 :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_1_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_1_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_1_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_1_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_1_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_1_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_1_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_1_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_1_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_1_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_1_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_1_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_1_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_1_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_1_upstream);
  --assign niosII_system_burst_1_upstream_readdata_from_sa = niosII_system_burst_1_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_1_upstream_readdata_from_sa <= niosII_system_burst_1_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_1_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("1100100001000100000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_1_upstream_waitrequest_from_sa = niosII_system_burst_1_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_1_upstream_waitrequest_from_sa <= niosII_system_burst_1_upstream_waitrequest;
  --assign niosII_system_burst_1_upstream_readdatavalid_from_sa = niosII_system_burst_1_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_1_upstream_readdatavalid_from_sa <= niosII_system_burst_1_upstream_readdatavalid;
  --niosII_system_burst_1_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_1_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_1_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_1_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_1_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_1_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_1_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_1_upstream;
  --niosII_system_burst_1_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_1_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_1_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_1_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_1_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_1_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_1_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_1_upstream_allgrants <= niosII_system_burst_1_upstream_grant_vector;
  --niosII_system_burst_1_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_1_upstream_end_xfer <= NOT ((niosII_system_burst_1_upstream_waits_for_read OR niosII_system_burst_1_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_1_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_1_upstream <= niosII_system_burst_1_upstream_end_xfer AND (((NOT niosII_system_burst_1_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_1_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_1_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_1_upstream AND niosII_system_burst_1_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_1_upstream AND NOT niosII_system_burst_1_upstream_non_bursting_master_requests));
  --niosII_system_burst_1_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_1_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_1_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_1_upstream_arb_share_counter <= niosII_system_burst_1_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_1_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_1_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_1_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_1_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_1_upstream AND NOT niosII_system_burst_1_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_1_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_1_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_1/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_1_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_1_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_1_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_1_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_1/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_1_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_1_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_1_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_1_upstream <= internal_cpu_data_master_requests_niosII_system_burst_1_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_1_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_1_upstream_move_on_to_next_transaction <= niosII_system_burst_1_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_1_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_1_upstream, which is an e_mux
  niosII_system_burst_1_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_1_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_1_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_1_upstream : burstcount_fifo_for_niosII_system_burst_1_upstream_module
    port map(
      data_out => niosII_system_burst_1_upstream_transaction_burst_count,
      empty => niosII_system_burst_1_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input6,
      clk => clk,
      data_in => niosII_system_burst_1_upstream_selected_burstcount,
      read => niosII_system_burst_1_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input7,
      write => module_input8
    );

  module_input6 <= std_logic'('0');
  module_input7 <= std_logic'('0');
  module_input8 <= ((in_a_read_cycle AND NOT niosII_system_burst_1_upstream_waits_for_read) AND niosII_system_burst_1_upstream_load_fifo) AND NOT ((niosII_system_burst_1_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_1_upstream_burstcount_fifo_empty));

  --niosII_system_burst_1_upstream current burst minus one, which is an e_assign
  niosII_system_burst_1_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_1_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_1_upstream, which is an e_mux
  niosII_system_burst_1_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_1_upstream_waits_for_read)) AND NOT niosII_system_burst_1_upstream_load_fifo))) = '1'), niosII_system_burst_1_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_1_upstream_waits_for_read) AND niosII_system_burst_1_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_1_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_1_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_1_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_1_upstream_transaction_burst_count, niosII_system_burst_1_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_1_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_1_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_1_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_1_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_1_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_1_upstream_current_burst <= niosII_system_burst_1_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_1_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_1_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_1_upstream_waits_for_read)) AND niosII_system_burst_1_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_1_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_1_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_1_upstream_waits_for_read)) AND NOT niosII_system_burst_1_upstream_load_fifo) OR niosII_system_burst_1_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_1_upstream_load_fifo <= p0_niosII_system_burst_1_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_1_upstream, which is an e_assign
  niosII_system_burst_1_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_1_upstream_current_burst_minus_one)) AND niosII_system_burst_1_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_1_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_1_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_1_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_1_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_1_upstream,
      full => open,
      clear_fifo => module_input9,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_1_upstream,
      read => niosII_system_burst_1_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input10,
      write => module_input11
    );

  module_input9 <= std_logic'('0');
  module_input10 <= std_logic'('0');
  module_input11 <= in_a_read_cycle AND NOT niosII_system_burst_1_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_1_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_1_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_1_upstream <= niosII_system_burst_1_upstream_readdatavalid_from_sa;
  --niosII_system_burst_1_upstream_writedata mux, which is an e_mux
  niosII_system_burst_1_upstream_writedata <= cpu_data_master_writedata;
  --byteaddress mux for niosII_system_burst_1/upstream, which is an e_mux
  niosII_system_burst_1_upstream_byteaddress <= cpu_data_master_address_to_slave (12 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_1_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_1_upstream;
  --cpu/data_master saved-grant niosII_system_burst_1/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_1_upstream <= internal_cpu_data_master_requests_niosII_system_burst_1_upstream;
  --allow new arb cycle for niosII_system_burst_1/upstream, which is an e_assign
  niosII_system_burst_1_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_1_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_1_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_1_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_1_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_1_upstream_begins_xfer) = '1'), niosII_system_burst_1_upstream_unreg_firsttransfer, niosII_system_burst_1_upstream_reg_firsttransfer);
  --niosII_system_burst_1_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_1_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_1_upstream_slavearbiterlockenable AND niosII_system_burst_1_upstream_any_continuerequest));
  --niosII_system_burst_1_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_1_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_1_upstream_begins_xfer) = '1' then 
        niosII_system_burst_1_upstream_reg_firsttransfer <= niosII_system_burst_1_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_1_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_1_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_1_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_1_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_1_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_1_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_1_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_1_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_1_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_1_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_1_upstream_begins_xfer) = '1' then 
        niosII_system_burst_1_upstream_bbt_burstcounter <= niosII_system_burst_1_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_1_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_1_upstream_beginbursttransfer_internal <= niosII_system_burst_1_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_1_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_1_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_1_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_1_upstream AND cpu_data_master_read;
  --niosII_system_burst_1_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_1_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_1_upstream AND cpu_data_master_write;
  --niosII_system_burst_1_upstream_address mux, which is an e_mux
  niosII_system_burst_1_upstream_address <= cpu_data_master_address_to_slave (10 DOWNTO 0);
  --d1_niosII_system_burst_1_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_1_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_1_upstream_end_xfer <= niosII_system_burst_1_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_1_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_1_upstream_waits_for_read <= niosII_system_burst_1_upstream_in_a_read_cycle AND internal_niosII_system_burst_1_upstream_waitrequest_from_sa;
  --niosII_system_burst_1_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_1_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_1_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_1_upstream_in_a_read_cycle;
  --niosII_system_burst_1_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_1_upstream_waits_for_write <= niosII_system_burst_1_upstream_in_a_write_cycle AND internal_niosII_system_burst_1_upstream_waitrequest_from_sa;
  --niosII_system_burst_1_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_1_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_1_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_1_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_1_upstream_counter <= std_logic'('0');
  --niosII_system_burst_1_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_1_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_1_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_1_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_1_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_1_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_1_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_1_upstream <= internal_cpu_data_master_granted_niosII_system_burst_1_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_1_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_1_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_1_upstream <= internal_cpu_data_master_requests_niosII_system_burst_1_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_1_upstream_burstcount <= internal_niosII_system_burst_1_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_1_upstream_read <= internal_niosII_system_burst_1_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_1_upstream_waitrequest_from_sa <= internal_niosII_system_burst_1_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_1_upstream_write <= internal_niosII_system_burst_1_upstream_write;
--synthesis translate_off
    --niosII_system_burst_1/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line38 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_1_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line38, now);
          write(write_line38, string'(": "));
          write(write_line38, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_1/upstream"));
          write(output, write_line38.all);
          deallocate (write_line38);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_1_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal niosII_system_burst_1_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_1_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal niosII_system_burst_1_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_1_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_1_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_1_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_1_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_1_downstream_arbitrator;


architecture europa of niosII_system_burst_1_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_1_downstream_address_to_slave :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal internal_niosII_system_burst_1_downstream_latency_counter :  STD_LOGIC;
                signal internal_niosII_system_burst_1_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_address_last_time :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_1_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_1_downstream_is_granted_some_slave :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_niosII_system_burst_1_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_niosII_system_burst_1_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module OR NOT niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module OR NOT niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module OR NOT niosII_system_burst_1_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cpu_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_1_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module OR NOT niosII_system_burst_1_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_1_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_1_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_1_downstream_address_to_slave <= niosII_system_burst_1_downstream_address;
  --niosII_system_burst_1_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_1_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_1_downstream_read_but_no_slave_selected <= (niosII_system_burst_1_downstream_read AND niosII_system_burst_1_downstream_run) AND NOT niosII_system_burst_1_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  niosII_system_burst_1_downstream_is_granted_some_slave <= niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_1_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_1_downstream_readdatavalid <= (niosII_system_burst_1_downstream_read_but_no_slave_selected OR pre_flush_niosII_system_burst_1_downstream_readdatavalid) OR niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module;
  --niosII_system_burst_1/downstream readdata mux, which is an e_mux
  niosII_system_burst_1_downstream_readdata <= cpu_jtag_debug_module_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_1_downstream_waitrequest <= NOT niosII_system_burst_1_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_niosII_system_burst_1_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_niosII_system_burst_1_downstream_latency_counter <= p1_niosII_system_burst_1_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_niosII_system_burst_1_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((niosII_system_burst_1_downstream_run AND niosII_system_burst_1_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_1_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_1_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --niosII_system_burst_1_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_1_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_1_downstream_address_to_slave <= internal_niosII_system_burst_1_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_1_downstream_latency_counter <= internal_niosII_system_burst_1_downstream_latency_counter;
  --vhdl renameroo for output signals
  niosII_system_burst_1_downstream_waitrequest <= internal_niosII_system_burst_1_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_1_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_1_downstream_address_last_time <= std_logic_vector'("00000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_1_downstream_address_last_time <= niosII_system_burst_1_downstream_address;
      end if;

    end process;

    --niosII_system_burst_1/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_1_downstream_waitrequest AND ((niosII_system_burst_1_downstream_read OR niosII_system_burst_1_downstream_write));
      end if;

    end process;

    --niosII_system_burst_1_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line39 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_1_downstream_address /= niosII_system_burst_1_downstream_address_last_time))))) = '1' then 
          write(write_line39, now);
          write(write_line39, string'(": "));
          write(write_line39, string'("niosII_system_burst_1_downstream_address did not heed wait!!!"));
          write(output, write_line39.all);
          deallocate (write_line39);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_1_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_1_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_1_downstream_burstcount_last_time <= niosII_system_burst_1_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_1_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line40 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_1_downstream_burstcount) /= std_logic'(niosII_system_burst_1_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line40, now);
          write(write_line40, string'(": "));
          write(write_line40, string'("niosII_system_burst_1_downstream_burstcount did not heed wait!!!"));
          write(output, write_line40.all);
          deallocate (write_line40);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_1_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_1_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_1_downstream_byteenable_last_time <= niosII_system_burst_1_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_1_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line41 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_1_downstream_byteenable /= niosII_system_burst_1_downstream_byteenable_last_time))))) = '1' then 
          write(write_line41, now);
          write(write_line41, string'(": "));
          write(write_line41, string'("niosII_system_burst_1_downstream_byteenable did not heed wait!!!"));
          write(output, write_line41.all);
          deallocate (write_line41);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_1_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_1_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_1_downstream_read_last_time <= niosII_system_burst_1_downstream_read;
      end if;

    end process;

    --niosII_system_burst_1_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line42 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_1_downstream_read) /= std_logic'(niosII_system_burst_1_downstream_read_last_time)))))) = '1' then 
          write(write_line42, now);
          write(write_line42, string'(": "));
          write(write_line42, string'("niosII_system_burst_1_downstream_read did not heed wait!!!"));
          write(output, write_line42.all);
          deallocate (write_line42);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_1_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_1_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_1_downstream_write_last_time <= niosII_system_burst_1_downstream_write;
      end if;

    end process;

    --niosII_system_burst_1_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line43 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_1_downstream_write) /= std_logic'(niosII_system_burst_1_downstream_write_last_time)))))) = '1' then 
          write(write_line43, now);
          write(write_line43, string'(": "));
          write(write_line43, string'("niosII_system_burst_1_downstream_write did not heed wait!!!"));
          write(output, write_line43.all);
          deallocate (write_line43);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_1_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_1_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_1_downstream_writedata_last_time <= niosII_system_burst_1_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_1_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line44 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_1_downstream_writedata /= niosII_system_burst_1_downstream_writedata_last_time)))) AND niosII_system_burst_1_downstream_write)) = '1' then 
          write(write_line44, now);
          write(write_line44, string'(": "));
          write(write_line44, string'("niosII_system_burst_1_downstream_writedata did not heed wait!!!"));
          write(output, write_line44.all);
          deallocate (write_line44);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_10_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_10_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_10_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_4 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_5 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_6 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_7 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_8 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic_vector'("00000");
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic_vector'("00000");
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic_vector'("00000");
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic_vector'("00000");
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic_vector'("00000");
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("00000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("00000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("00000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("00000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_10_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_10_upstream_module;


architecture europa of rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_10_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_10_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : IN STD_LOGIC;
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : IN STD_LOGIC;
                 signal niosII_system_burst_10_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_10_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_10_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_instruction_master_granted_niosII_system_burst_10_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_instruction_master_requests_niosII_system_burst_10_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_10_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_10_upstream_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal niosII_system_burst_10_upstream_byteaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal niosII_system_burst_10_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_10_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_10_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_10_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_10_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_10_upstream_write : OUT STD_LOGIC
              );
end entity niosII_system_burst_10_upstream_arbitrator;


architecture europa of niosII_system_burst_10_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_10_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_10_upstream_module;

component rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_10_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_10_upstream_module;

                signal cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_output_from_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal cpu_instruction_master_saved_grant_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_instruction_master_granted_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal internal_cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal internal_cpu_instruction_master_requests_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_10_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal module_input12 :  STD_LOGIC;
                signal module_input13 :  STD_LOGIC;
                signal module_input14 :  STD_LOGIC;
                signal module_input15 :  STD_LOGIC;
                signal module_input16 :  STD_LOGIC;
                signal module_input17 :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_10_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_10_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_10_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_current_burst :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_10_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_10_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_next_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_10_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_selected_burstcount :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_10_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_10_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_10_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_10_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_10_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_10_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream);
  --assign niosII_system_burst_10_upstream_readdatavalid_from_sa = niosII_system_burst_10_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_10_upstream_readdatavalid_from_sa <= niosII_system_burst_10_upstream_readdatavalid;
  --assign niosII_system_burst_10_upstream_readdata_from_sa = niosII_system_burst_10_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_10_upstream_readdata_from_sa <= niosII_system_burst_10_upstream_readdata;
  internal_cpu_instruction_master_requests_niosII_system_burst_10_upstream <= ((to_std_logic(((Std_Logic_Vector'(cpu_instruction_master_address_to_slave(24 DOWNTO 23) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("0100000000000000000000000")))) AND (cpu_instruction_master_read))) AND cpu_instruction_master_read;
  --assign niosII_system_burst_10_upstream_waitrequest_from_sa = niosII_system_burst_10_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_10_upstream_waitrequest_from_sa <= niosII_system_burst_10_upstream_waitrequest;
  --niosII_system_burst_10_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_10_upstream_arb_share_set_values <= std_logic_vector'("00000001");
  --niosII_system_burst_10_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_10_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_10_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_10_upstream_any_bursting_master_saved_grant <= cpu_instruction_master_saved_grant_niosII_system_burst_10_upstream;
  --niosII_system_burst_10_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_10_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_10_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_10_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_10_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_10_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_10_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_10_upstream_allgrants <= niosII_system_burst_10_upstream_grant_vector;
  --niosII_system_burst_10_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_10_upstream_end_xfer <= NOT ((niosII_system_burst_10_upstream_waits_for_read OR niosII_system_burst_10_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_10_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_10_upstream <= niosII_system_burst_10_upstream_end_xfer AND (((NOT niosII_system_burst_10_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_10_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_10_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_10_upstream AND niosII_system_burst_10_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_10_upstream AND NOT niosII_system_burst_10_upstream_non_bursting_master_requests));
  --niosII_system_burst_10_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_10_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_10_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_10_upstream_arb_share_counter <= niosII_system_burst_10_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_10_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_10_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_10_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_10_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_10_upstream AND NOT niosII_system_burst_10_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_10_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_10_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/instruction_master niosII_system_burst_10/upstream arbiterlock, which is an e_assign
  cpu_instruction_master_arbiterlock <= niosII_system_burst_10_upstream_slavearbiterlockenable AND cpu_instruction_master_continuerequest;
  --niosII_system_burst_10_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_10_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_10_upstream_arb_share_counter_next_value);
  --cpu/instruction_master niosII_system_burst_10/upstream arbiterlock2, which is an e_assign
  cpu_instruction_master_arbiterlock2 <= niosII_system_burst_10_upstream_slavearbiterlockenable2 AND cpu_instruction_master_continuerequest;
  --niosII_system_burst_10_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_10_upstream_any_continuerequest <= std_logic'('1');
  --cpu_instruction_master_continuerequest continued request, which is an e_assign
  cpu_instruction_master_continuerequest <= std_logic'('1');
  internal_cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_10_upstream AND NOT ((cpu_instruction_master_read AND (((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_latency_counter))))))) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register)))));
  --unique name for niosII_system_burst_10_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_10_upstream_move_on_to_next_transaction <= niosII_system_burst_10_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_10_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_10_upstream, which is an e_mux
  niosII_system_burst_10_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_niosII_system_burst_10_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_instruction_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --burstcount_fifo_for_niosII_system_burst_10_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_10_upstream : burstcount_fifo_for_niosII_system_burst_10_upstream_module
    port map(
      data_out => niosII_system_burst_10_upstream_transaction_burst_count,
      empty => niosII_system_burst_10_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input12,
      clk => clk,
      data_in => niosII_system_burst_10_upstream_selected_burstcount,
      read => niosII_system_burst_10_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input13,
      write => module_input14
    );

  module_input12 <= std_logic'('0');
  module_input13 <= std_logic'('0');
  module_input14 <= ((in_a_read_cycle AND NOT niosII_system_burst_10_upstream_waits_for_read) AND niosII_system_burst_10_upstream_load_fifo) AND NOT ((niosII_system_burst_10_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_10_upstream_burstcount_fifo_empty));

  --niosII_system_burst_10_upstream current burst minus one, which is an e_assign
  niosII_system_burst_10_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_10_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --what to load in current_burst, for niosII_system_burst_10_upstream, which is an e_mux
  niosII_system_burst_10_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_10_upstream_waits_for_read)) AND NOT niosII_system_burst_10_upstream_load_fifo))) = '1'), (niosII_system_burst_10_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_10_upstream_waits_for_read) AND niosII_system_burst_10_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_10_upstream_burstcount_fifo_empty))) = '1'), (niosII_system_burst_10_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'((niosII_system_burst_10_upstream_this_cycle_is_the_last_burst)) = '1'), (niosII_system_burst_10_upstream_transaction_burst_count & A_ToStdLogicVector(std_logic'('0'))), (std_logic_vector'("0") & (niosII_system_burst_10_upstream_current_burst_minus_one))))), 5);
  --the current burst count for niosII_system_burst_10_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_10_upstream_current_burst <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_10_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_10_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_10_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_10_upstream_current_burst <= niosII_system_burst_10_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_10_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_10_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_10_upstream_waits_for_read)) AND niosII_system_burst_10_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_10_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_10_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_10_upstream_waits_for_read)) AND NOT niosII_system_burst_10_upstream_load_fifo) OR niosII_system_burst_10_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_10_upstream_load_fifo <= p0_niosII_system_burst_10_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_10_upstream, which is an e_assign
  niosII_system_burst_10_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_10_upstream_current_burst_minus_one)) AND niosII_system_burst_10_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_10_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_10_upstream : rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_10_upstream_module
    port map(
      data_out => cpu_instruction_master_rdv_fifo_output_from_niosII_system_burst_10_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_10_upstream,
      full => open,
      clear_fifo => module_input15,
      clk => clk,
      data_in => internal_cpu_instruction_master_granted_niosII_system_burst_10_upstream,
      read => niosII_system_burst_10_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input16,
      write => module_input17
    );

  module_input15 <= std_logic'('0');
  module_input16 <= std_logic'('0');
  module_input17 <= in_a_read_cycle AND NOT niosII_system_burst_10_upstream_waits_for_read;

  cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register <= NOT cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_10_upstream;
  --local readdatavalid cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream, which is an e_mux
  cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream <= niosII_system_burst_10_upstream_readdatavalid_from_sa;
  --byteaddress mux for niosII_system_burst_10/upstream, which is an e_mux
  niosII_system_burst_10_upstream_byteaddress <= cpu_instruction_master_address_to_slave (23 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_instruction_master_granted_niosII_system_burst_10_upstream <= internal_cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream;
  --cpu/instruction_master saved-grant niosII_system_burst_10/upstream, which is an e_assign
  cpu_instruction_master_saved_grant_niosII_system_burst_10_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_10_upstream;
  --allow new arb cycle for niosII_system_burst_10/upstream, which is an e_assign
  niosII_system_burst_10_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_10_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_10_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_10_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_10_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_10_upstream_begins_xfer) = '1'), niosII_system_burst_10_upstream_unreg_firsttransfer, niosII_system_burst_10_upstream_reg_firsttransfer);
  --niosII_system_burst_10_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_10_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_10_upstream_slavearbiterlockenable AND niosII_system_burst_10_upstream_any_continuerequest));
  --niosII_system_burst_10_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_10_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_10_upstream_begins_xfer) = '1' then 
        niosII_system_burst_10_upstream_reg_firsttransfer <= niosII_system_burst_10_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_10_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_10_upstream_beginbursttransfer_internal <= niosII_system_burst_10_upstream_begins_xfer;
  --niosII_system_burst_10_upstream_read assignment, which is an e_mux
  niosII_system_burst_10_upstream_read <= internal_cpu_instruction_master_granted_niosII_system_burst_10_upstream AND cpu_instruction_master_read;
  --niosII_system_burst_10_upstream_write assignment, which is an e_mux
  niosII_system_burst_10_upstream_write <= std_logic'('0');
  --niosII_system_burst_10_upstream_address mux, which is an e_mux
  niosII_system_burst_10_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(cpu_instruction_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 23);
  --d1_niosII_system_burst_10_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_10_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_10_upstream_end_xfer <= niosII_system_burst_10_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_10_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_10_upstream_waits_for_read <= niosII_system_burst_10_upstream_in_a_read_cycle AND internal_niosII_system_burst_10_upstream_waitrequest_from_sa;
  --niosII_system_burst_10_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_10_upstream_in_a_read_cycle <= internal_cpu_instruction_master_granted_niosII_system_burst_10_upstream AND cpu_instruction_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_10_upstream_in_a_read_cycle;
  --niosII_system_burst_10_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_10_upstream_waits_for_write <= niosII_system_burst_10_upstream_in_a_write_cycle AND internal_niosII_system_burst_10_upstream_waitrequest_from_sa;
  --niosII_system_burst_10_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_10_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_10_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_10_upstream_counter <= std_logic'('0');
  --niosII_system_burst_10_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_10_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 2);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_10_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_instruction_master_granted_niosII_system_burst_10_upstream <= internal_cpu_instruction_master_granted_niosII_system_burst_10_upstream;
  --vhdl renameroo for output signals
  cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream <= internal_cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream;
  --vhdl renameroo for output signals
  cpu_instruction_master_requests_niosII_system_burst_10_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_10_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_10_upstream_waitrequest_from_sa <= internal_niosII_system_burst_10_upstream_waitrequest_from_sa;
--synthesis translate_off
    --niosII_system_burst_10/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/instruction_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line45 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_instruction_master_requests_niosII_system_burst_10_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_instruction_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line45, now);
          write(write_line45, string'(": "));
          write(write_line45, string'("cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_10/upstream"));
          write(output, write_line45.all);
          deallocate (write_line45);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_10_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal niosII_system_burst_10_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_10_downstream_granted_sdram_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_requests_sdram_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_10_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal niosII_system_burst_10_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_10_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_10_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_10_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_10_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_10_downstream_arbitrator;


architecture europa of niosII_system_burst_10_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_10_downstream_address_to_slave :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal internal_niosII_system_burst_10_downstream_latency_counter :  STD_LOGIC;
                signal internal_niosII_system_burst_10_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_address_last_time :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_10_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_10_downstream_is_granted_some_slave :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_niosII_system_burst_10_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_niosII_system_burst_10_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_10_downstream_qualified_request_sdram_s1 OR NOT niosII_system_burst_10_downstream_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_10_downstream_granted_sdram_s1 OR NOT niosII_system_burst_10_downstream_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_10_downstream_qualified_request_sdram_s1 OR NOT ((niosII_system_burst_10_downstream_read OR niosII_system_burst_10_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_10_downstream_read OR niosII_system_burst_10_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_10_downstream_qualified_request_sdram_s1 OR NOT ((niosII_system_burst_10_downstream_read OR niosII_system_burst_10_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_10_downstream_read OR niosII_system_burst_10_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_10_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_10_downstream_address_to_slave <= niosII_system_burst_10_downstream_address;
  --niosII_system_burst_10_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_10_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_10_downstream_read_but_no_slave_selected <= (niosII_system_burst_10_downstream_read AND niosII_system_burst_10_downstream_run) AND NOT niosII_system_burst_10_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  niosII_system_burst_10_downstream_is_granted_some_slave <= niosII_system_burst_10_downstream_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_10_downstream_readdatavalid <= niosII_system_burst_10_downstream_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_10_downstream_readdatavalid <= niosII_system_burst_10_downstream_read_but_no_slave_selected OR pre_flush_niosII_system_burst_10_downstream_readdatavalid;
  --niosII_system_burst_10/downstream readdata mux, which is an e_mux
  niosII_system_burst_10_downstream_readdata <= sdram_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_10_downstream_waitrequest <= NOT niosII_system_burst_10_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_niosII_system_burst_10_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_niosII_system_burst_10_downstream_latency_counter <= p1_niosII_system_burst_10_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_niosII_system_burst_10_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((niosII_system_burst_10_downstream_run AND niosII_system_burst_10_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_10_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_10_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --niosII_system_burst_10_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_10_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_10_downstream_address_to_slave <= internal_niosII_system_burst_10_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_10_downstream_latency_counter <= internal_niosII_system_burst_10_downstream_latency_counter;
  --vhdl renameroo for output signals
  niosII_system_burst_10_downstream_waitrequest <= internal_niosII_system_burst_10_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_10_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_10_downstream_address_last_time <= std_logic_vector'("00000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_10_downstream_address_last_time <= niosII_system_burst_10_downstream_address;
      end if;

    end process;

    --niosII_system_burst_10/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_10_downstream_waitrequest AND ((niosII_system_burst_10_downstream_read OR niosII_system_burst_10_downstream_write));
      end if;

    end process;

    --niosII_system_burst_10_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line46 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_10_downstream_address /= niosII_system_burst_10_downstream_address_last_time))))) = '1' then 
          write(write_line46, now);
          write(write_line46, string'(": "));
          write(write_line46, string'("niosII_system_burst_10_downstream_address did not heed wait!!!"));
          write(output, write_line46.all);
          deallocate (write_line46);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_10_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_10_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_10_downstream_burstcount_last_time <= niosII_system_burst_10_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_10_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line47 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_10_downstream_burstcount) /= std_logic'(niosII_system_burst_10_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line47, now);
          write(write_line47, string'(": "));
          write(write_line47, string'("niosII_system_burst_10_downstream_burstcount did not heed wait!!!"));
          write(output, write_line47.all);
          deallocate (write_line47);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_10_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_10_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_10_downstream_byteenable_last_time <= niosII_system_burst_10_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_10_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line48 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_10_downstream_byteenable /= niosII_system_burst_10_downstream_byteenable_last_time))))) = '1' then 
          write(write_line48, now);
          write(write_line48, string'(": "));
          write(write_line48, string'("niosII_system_burst_10_downstream_byteenable did not heed wait!!!"));
          write(output, write_line48.all);
          deallocate (write_line48);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_10_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_10_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_10_downstream_read_last_time <= niosII_system_burst_10_downstream_read;
      end if;

    end process;

    --niosII_system_burst_10_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line49 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_10_downstream_read) /= std_logic'(niosII_system_burst_10_downstream_read_last_time)))))) = '1' then 
          write(write_line49, now);
          write(write_line49, string'(": "));
          write(write_line49, string'("niosII_system_burst_10_downstream_read did not heed wait!!!"));
          write(output, write_line49.all);
          deallocate (write_line49);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_10_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_10_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_10_downstream_write_last_time <= niosII_system_burst_10_downstream_write;
      end if;

    end process;

    --niosII_system_burst_10_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line50 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_10_downstream_write) /= std_logic'(niosII_system_burst_10_downstream_write_last_time)))))) = '1' then 
          write(write_line50, now);
          write(write_line50, string'(": "));
          write(write_line50, string'("niosII_system_burst_10_downstream_write did not heed wait!!!"));
          write(output, write_line50.all);
          deallocate (write_line50);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_10_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_10_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_10_downstream_writedata_last_time <= niosII_system_burst_10_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_10_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line51 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_10_downstream_writedata /= niosII_system_burst_10_downstream_writedata_last_time)))) AND niosII_system_burst_10_downstream_write)) = '1' then 
          write(write_line51, now);
          write(write_line51, string'(": "));
          write(write_line51, string'("niosII_system_burst_10_downstream_writedata did not heed wait!!!"));
          write(output, write_line51.all);
          deallocate (write_line51);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_11_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_11_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_11_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_4 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_5 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_6 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_7 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_8 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic_vector'("00000");
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic_vector'("00000");
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic_vector'("00000");
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic_vector'("00000");
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic_vector'("00000");
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("00000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("00000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("00000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("00000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_11_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_11_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_11_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_11_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal niosII_system_burst_11_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_11_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_11_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_byteenable_niosII_system_burst_11_upstream : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_granted_niosII_system_burst_11_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_11_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_11_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_11_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_11_upstream_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal niosII_system_burst_11_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_11_upstream_byteaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal niosII_system_burst_11_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_11_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_11_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_11_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_11_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_11_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_11_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity niosII_system_burst_11_upstream_arbitrator;


architecture europa of niosII_system_burst_11_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_11_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_11_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_11_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_11_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_byteenable_niosII_system_burst_11_upstream_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_byteenable_niosII_system_burst_11_upstream_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_byteenable_niosII_system_burst_11_upstream :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_data_master_granted_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_11_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_11_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_11_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_11_upstream_write :  STD_LOGIC;
                signal module_input18 :  STD_LOGIC;
                signal module_input19 :  STD_LOGIC;
                signal module_input20 :  STD_LOGIC;
                signal module_input21 :  STD_LOGIC;
                signal module_input22 :  STD_LOGIC;
                signal module_input23 :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_11_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_11_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_11_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_11_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_current_burst :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_11_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_11_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_11_upstream_next_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_11_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_selected_burstcount :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_11_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_11_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_11_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_11_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_11_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_11_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_11_upstream);
  --assign niosII_system_burst_11_upstream_readdatavalid_from_sa = niosII_system_burst_11_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_11_upstream_readdatavalid_from_sa <= niosII_system_burst_11_upstream_readdatavalid;
  --assign niosII_system_burst_11_upstream_readdata_from_sa = niosII_system_burst_11_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_11_upstream_readdata_from_sa <= niosII_system_burst_11_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_11_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 23) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("0100000000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_11_upstream_waitrequest_from_sa = niosII_system_burst_11_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_11_upstream_waitrequest_from_sa <= niosII_system_burst_11_upstream_waitrequest;
  --niosII_system_burst_11_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_11_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_11_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (A_SLL(cpu_data_master_burstcount,std_logic_vector'("00000000000000000000000000000001")))), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_11_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_11_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_11_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_11_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_11_upstream;
  --niosII_system_burst_11_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_11_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_11_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_11_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_11_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_11_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_11_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_11_upstream_allgrants <= niosII_system_burst_11_upstream_grant_vector;
  --niosII_system_burst_11_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_11_upstream_end_xfer <= NOT ((niosII_system_burst_11_upstream_waits_for_read OR niosII_system_burst_11_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_11_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_11_upstream <= niosII_system_burst_11_upstream_end_xfer AND (((NOT niosII_system_burst_11_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_11_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_11_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_11_upstream AND niosII_system_burst_11_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_11_upstream AND NOT niosII_system_burst_11_upstream_non_bursting_master_requests));
  --niosII_system_burst_11_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_11_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_11_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_11_upstream_arb_share_counter <= niosII_system_burst_11_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_11_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_11_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_11_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_11_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_11_upstream AND NOT niosII_system_burst_11_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_11_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_11_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_11/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_11_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_11_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_11_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_11_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_11/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_11_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_11_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_11_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_11_upstream <= internal_cpu_data_master_requests_niosII_system_burst_11_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_11_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_11_upstream_move_on_to_next_transaction <= niosII_system_burst_11_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_11_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_11_upstream, which is an e_mux
  niosII_system_burst_11_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_11_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --burstcount_fifo_for_niosII_system_burst_11_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_11_upstream : burstcount_fifo_for_niosII_system_burst_11_upstream_module
    port map(
      data_out => niosII_system_burst_11_upstream_transaction_burst_count,
      empty => niosII_system_burst_11_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input18,
      clk => clk,
      data_in => niosII_system_burst_11_upstream_selected_burstcount,
      read => niosII_system_burst_11_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input19,
      write => module_input20
    );

  module_input18 <= std_logic'('0');
  module_input19 <= std_logic'('0');
  module_input20 <= ((in_a_read_cycle AND NOT niosII_system_burst_11_upstream_waits_for_read) AND niosII_system_burst_11_upstream_load_fifo) AND NOT ((niosII_system_burst_11_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_11_upstream_burstcount_fifo_empty));

  --niosII_system_burst_11_upstream current burst minus one, which is an e_assign
  niosII_system_burst_11_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_11_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --what to load in current_burst, for niosII_system_burst_11_upstream, which is an e_mux
  niosII_system_burst_11_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_11_upstream_waits_for_read)) AND NOT niosII_system_burst_11_upstream_load_fifo))) = '1'), (niosII_system_burst_11_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_11_upstream_waits_for_read) AND niosII_system_burst_11_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_11_upstream_burstcount_fifo_empty))) = '1'), (niosII_system_burst_11_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'((niosII_system_burst_11_upstream_this_cycle_is_the_last_burst)) = '1'), (niosII_system_burst_11_upstream_transaction_burst_count & A_ToStdLogicVector(std_logic'('0'))), (std_logic_vector'("0") & (niosII_system_burst_11_upstream_current_burst_minus_one))))), 5);
  --the current burst count for niosII_system_burst_11_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_11_upstream_current_burst <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_11_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_11_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_11_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_11_upstream_current_burst <= niosII_system_burst_11_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_11_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_11_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_11_upstream_waits_for_read)) AND niosII_system_burst_11_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_11_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_11_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_11_upstream_waits_for_read)) AND NOT niosII_system_burst_11_upstream_load_fifo) OR niosII_system_burst_11_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_11_upstream_load_fifo <= p0_niosII_system_burst_11_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_11_upstream, which is an e_assign
  niosII_system_burst_11_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_11_upstream_current_burst_minus_one)) AND niosII_system_burst_11_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_11_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_11_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_11_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_11_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_11_upstream,
      full => open,
      clear_fifo => module_input21,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_11_upstream,
      read => niosII_system_burst_11_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input22,
      write => module_input23
    );

  module_input21 <= std_logic'('0');
  module_input22 <= std_logic'('0');
  module_input23 <= in_a_read_cycle AND NOT niosII_system_burst_11_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_11_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_11_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_11_upstream <= niosII_system_burst_11_upstream_readdatavalid_from_sa;
  --niosII_system_burst_11_upstream_writedata mux, which is an e_mux
  niosII_system_burst_11_upstream_writedata <= cpu_data_master_dbs_write_16;
  --byteaddress mux for niosII_system_burst_11/upstream, which is an e_mux
  niosII_system_burst_11_upstream_byteaddress <= cpu_data_master_address_to_slave (23 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_11_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_11_upstream;
  --cpu/data_master saved-grant niosII_system_burst_11/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_11_upstream <= internal_cpu_data_master_requests_niosII_system_burst_11_upstream;
  --allow new arb cycle for niosII_system_burst_11/upstream, which is an e_assign
  niosII_system_burst_11_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_11_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_11_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_11_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_11_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_11_upstream_begins_xfer) = '1'), niosII_system_burst_11_upstream_unreg_firsttransfer, niosII_system_burst_11_upstream_reg_firsttransfer);
  --niosII_system_burst_11_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_11_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_11_upstream_slavearbiterlockenable AND niosII_system_burst_11_upstream_any_continuerequest));
  --niosII_system_burst_11_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_11_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_11_upstream_begins_xfer) = '1' then 
        niosII_system_burst_11_upstream_reg_firsttransfer <= niosII_system_burst_11_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_11_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_11_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_11_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_11_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_11_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_11_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_11_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_11_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_11_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_11_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_11_upstream_begins_xfer) = '1' then 
        niosII_system_burst_11_upstream_bbt_burstcounter <= niosII_system_burst_11_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_11_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_11_upstream_beginbursttransfer_internal <= niosII_system_burst_11_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_11_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_11_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_11_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_11_upstream AND cpu_data_master_read;
  --niosII_system_burst_11_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_11_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_11_upstream AND cpu_data_master_write;
  --niosII_system_burst_11_upstream_address mux, which is an e_mux
  niosII_system_burst_11_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(cpu_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 23);
  --d1_niosII_system_burst_11_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_11_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_11_upstream_end_xfer <= niosII_system_burst_11_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_11_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_11_upstream_waits_for_read <= niosII_system_burst_11_upstream_in_a_read_cycle AND internal_niosII_system_burst_11_upstream_waitrequest_from_sa;
  --niosII_system_burst_11_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_11_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_11_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_11_upstream_in_a_read_cycle;
  --niosII_system_burst_11_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_11_upstream_waits_for_write <= niosII_system_burst_11_upstream_in_a_write_cycle AND internal_niosII_system_burst_11_upstream_waitrequest_from_sa;
  --niosII_system_burst_11_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_11_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_11_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_11_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_11_upstream_counter <= std_logic'('0');
  --niosII_system_burst_11_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_11_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_11_upstream)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_byteenable_niosII_system_burst_11_upstream)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  (cpu_data_master_byteenable_niosII_system_burst_11_upstream_segment_1(1), cpu_data_master_byteenable_niosII_system_burst_11_upstream_segment_1(0), cpu_data_master_byteenable_niosII_system_burst_11_upstream_segment_0(1), cpu_data_master_byteenable_niosII_system_burst_11_upstream_segment_0(0)) <= cpu_data_master_byteenable;
  internal_cpu_data_master_byteenable_niosII_system_burst_11_upstream <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), cpu_data_master_byteenable_niosII_system_burst_11_upstream_segment_0, cpu_data_master_byteenable_niosII_system_burst_11_upstream_segment_1);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_11_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_11_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_11_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_11_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_byteenable_niosII_system_burst_11_upstream <= internal_cpu_data_master_byteenable_niosII_system_burst_11_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_11_upstream <= internal_cpu_data_master_granted_niosII_system_burst_11_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_11_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_11_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_11_upstream <= internal_cpu_data_master_requests_niosII_system_burst_11_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_11_upstream_burstcount <= internal_niosII_system_burst_11_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_11_upstream_read <= internal_niosII_system_burst_11_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_11_upstream_waitrequest_from_sa <= internal_niosII_system_burst_11_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_11_upstream_write <= internal_niosII_system_burst_11_upstream_write;
--synthesis translate_off
    --niosII_system_burst_11/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line52 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_11_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line52, now);
          write(write_line52, string'(": "));
          write(write_line52, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_11/upstream"));
          write(output, write_line52.all);
          deallocate (write_line52);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_11_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal niosII_system_burst_11_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_11_downstream_granted_sdram_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_requests_sdram_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_11_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal niosII_system_burst_11_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_11_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_11_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_11_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_11_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_11_downstream_arbitrator;


architecture europa of niosII_system_burst_11_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_11_downstream_address_to_slave :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal internal_niosII_system_burst_11_downstream_latency_counter :  STD_LOGIC;
                signal internal_niosII_system_burst_11_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_address_last_time :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_11_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_11_downstream_is_granted_some_slave :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_niosII_system_burst_11_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_niosII_system_burst_11_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_11_downstream_qualified_request_sdram_s1 OR NOT niosII_system_burst_11_downstream_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_11_downstream_granted_sdram_s1 OR NOT niosII_system_burst_11_downstream_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_11_downstream_qualified_request_sdram_s1 OR NOT ((niosII_system_burst_11_downstream_read OR niosII_system_burst_11_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_11_downstream_read OR niosII_system_burst_11_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_11_downstream_qualified_request_sdram_s1 OR NOT ((niosII_system_burst_11_downstream_read OR niosII_system_burst_11_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_11_downstream_read OR niosII_system_burst_11_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_11_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_11_downstream_address_to_slave <= niosII_system_burst_11_downstream_address;
  --niosII_system_burst_11_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_11_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_11_downstream_read_but_no_slave_selected <= (niosII_system_burst_11_downstream_read AND niosII_system_burst_11_downstream_run) AND NOT niosII_system_burst_11_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  niosII_system_burst_11_downstream_is_granted_some_slave <= niosII_system_burst_11_downstream_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_11_downstream_readdatavalid <= niosII_system_burst_11_downstream_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_11_downstream_readdatavalid <= niosII_system_burst_11_downstream_read_but_no_slave_selected OR pre_flush_niosII_system_burst_11_downstream_readdatavalid;
  --niosII_system_burst_11/downstream readdata mux, which is an e_mux
  niosII_system_burst_11_downstream_readdata <= sdram_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_11_downstream_waitrequest <= NOT niosII_system_burst_11_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_niosII_system_burst_11_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_niosII_system_burst_11_downstream_latency_counter <= p1_niosII_system_burst_11_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_niosII_system_burst_11_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((niosII_system_burst_11_downstream_run AND niosII_system_burst_11_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_11_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_11_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --niosII_system_burst_11_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_11_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_11_downstream_address_to_slave <= internal_niosII_system_burst_11_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_11_downstream_latency_counter <= internal_niosII_system_burst_11_downstream_latency_counter;
  --vhdl renameroo for output signals
  niosII_system_burst_11_downstream_waitrequest <= internal_niosII_system_burst_11_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_11_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_11_downstream_address_last_time <= std_logic_vector'("00000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_11_downstream_address_last_time <= niosII_system_burst_11_downstream_address;
      end if;

    end process;

    --niosII_system_burst_11/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_11_downstream_waitrequest AND ((niosII_system_burst_11_downstream_read OR niosII_system_burst_11_downstream_write));
      end if;

    end process;

    --niosII_system_burst_11_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line53 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_11_downstream_address /= niosII_system_burst_11_downstream_address_last_time))))) = '1' then 
          write(write_line53, now);
          write(write_line53, string'(": "));
          write(write_line53, string'("niosII_system_burst_11_downstream_address did not heed wait!!!"));
          write(output, write_line53.all);
          deallocate (write_line53);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_11_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_11_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_11_downstream_burstcount_last_time <= niosII_system_burst_11_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_11_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line54 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_11_downstream_burstcount) /= std_logic'(niosII_system_burst_11_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line54, now);
          write(write_line54, string'(": "));
          write(write_line54, string'("niosII_system_burst_11_downstream_burstcount did not heed wait!!!"));
          write(output, write_line54.all);
          deallocate (write_line54);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_11_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_11_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_11_downstream_byteenable_last_time <= niosII_system_burst_11_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_11_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line55 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_11_downstream_byteenable /= niosII_system_burst_11_downstream_byteenable_last_time))))) = '1' then 
          write(write_line55, now);
          write(write_line55, string'(": "));
          write(write_line55, string'("niosII_system_burst_11_downstream_byteenable did not heed wait!!!"));
          write(output, write_line55.all);
          deallocate (write_line55);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_11_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_11_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_11_downstream_read_last_time <= niosII_system_burst_11_downstream_read;
      end if;

    end process;

    --niosII_system_burst_11_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line56 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_11_downstream_read) /= std_logic'(niosII_system_burst_11_downstream_read_last_time)))))) = '1' then 
          write(write_line56, now);
          write(write_line56, string'(": "));
          write(write_line56, string'("niosII_system_burst_11_downstream_read did not heed wait!!!"));
          write(output, write_line56.all);
          deallocate (write_line56);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_11_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_11_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_11_downstream_write_last_time <= niosII_system_burst_11_downstream_write;
      end if;

    end process;

    --niosII_system_burst_11_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line57 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_11_downstream_write) /= std_logic'(niosII_system_burst_11_downstream_write_last_time)))))) = '1' then 
          write(write_line57, now);
          write(write_line57, string'(": "));
          write(write_line57, string'("niosII_system_burst_11_downstream_write did not heed wait!!!"));
          write(output, write_line57.all);
          deallocate (write_line57);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_11_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_11_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_11_downstream_writedata_last_time <= niosII_system_burst_11_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_11_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line58 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_11_downstream_writedata /= niosII_system_burst_11_downstream_writedata_last_time)))) AND niosII_system_burst_11_downstream_write)) = '1' then 
          write(write_line58, now);
          write(write_line58, string'(": "));
          write(write_line58, string'("niosII_system_burst_11_downstream_writedata did not heed wait!!!"));
          write(output, write_line58.all);
          deallocate (write_line58);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_12_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_12_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_12_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("000000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("000000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("000000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("000000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_12_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_12_upstream_module;


architecture europa of rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_12_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_12_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : IN STD_LOGIC;
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : IN STD_LOGIC;
                 signal niosII_system_burst_12_upstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_12_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_12_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_instruction_master_granted_niosII_system_burst_12_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_instruction_master_requests_niosII_system_burst_12_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_12_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_12_upstream_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal niosII_system_burst_12_upstream_byteaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal niosII_system_burst_12_upstream_byteenable : OUT STD_LOGIC;
                 signal niosII_system_burst_12_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_12_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_12_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_12_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_12_upstream_write : OUT STD_LOGIC
              );
end entity niosII_system_burst_12_upstream_arbitrator;


architecture europa of niosII_system_burst_12_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_12_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_12_upstream_module;

component rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_12_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_12_upstream_module;

                signal cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_output_from_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal cpu_instruction_master_saved_grant_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_instruction_master_granted_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal internal_cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal internal_cpu_instruction_master_requests_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_12_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal module_input24 :  STD_LOGIC;
                signal module_input25 :  STD_LOGIC;
                signal module_input26 :  STD_LOGIC;
                signal module_input27 :  STD_LOGIC;
                signal module_input28 :  STD_LOGIC;
                signal module_input29 :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_12_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_12_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_12_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_current_burst :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_12_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_12_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_next_burst_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_12_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_selected_burstcount :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_12_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_12_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_12_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_12_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_12_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_12_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream);
  --assign niosII_system_burst_12_upstream_readdatavalid_from_sa = niosII_system_burst_12_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_12_upstream_readdatavalid_from_sa <= niosII_system_burst_12_upstream_readdatavalid;
  --assign niosII_system_burst_12_upstream_readdata_from_sa = niosII_system_burst_12_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_12_upstream_readdata_from_sa <= niosII_system_burst_12_upstream_readdata;
  internal_cpu_instruction_master_requests_niosII_system_burst_12_upstream <= ((to_std_logic(((Std_Logic_Vector'(cpu_instruction_master_address_to_slave(24 DOWNTO 22) & std_logic_vector'("0000000000000000000000")) = std_logic_vector'("1010000000000000000000000")))) AND (cpu_instruction_master_read))) AND cpu_instruction_master_read;
  --assign niosII_system_burst_12_upstream_waitrequest_from_sa = niosII_system_burst_12_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_12_upstream_waitrequest_from_sa <= niosII_system_burst_12_upstream_waitrequest;
  --niosII_system_burst_12_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_12_upstream_arb_share_set_values <= std_logic_vector'("00000001");
  --niosII_system_burst_12_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_12_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_12_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_12_upstream_any_bursting_master_saved_grant <= cpu_instruction_master_saved_grant_niosII_system_burst_12_upstream;
  --niosII_system_burst_12_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_12_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_12_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_12_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_12_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_12_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_12_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_12_upstream_allgrants <= niosII_system_burst_12_upstream_grant_vector;
  --niosII_system_burst_12_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_12_upstream_end_xfer <= NOT ((niosII_system_burst_12_upstream_waits_for_read OR niosII_system_burst_12_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_12_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_12_upstream <= niosII_system_burst_12_upstream_end_xfer AND (((NOT niosII_system_burst_12_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_12_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_12_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_12_upstream AND niosII_system_burst_12_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_12_upstream AND NOT niosII_system_burst_12_upstream_non_bursting_master_requests));
  --niosII_system_burst_12_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_12_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_12_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_12_upstream_arb_share_counter <= niosII_system_burst_12_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_12_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_12_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_12_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_12_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_12_upstream AND NOT niosII_system_burst_12_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_12_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_12_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/instruction_master niosII_system_burst_12/upstream arbiterlock, which is an e_assign
  cpu_instruction_master_arbiterlock <= niosII_system_burst_12_upstream_slavearbiterlockenable AND cpu_instruction_master_continuerequest;
  --niosII_system_burst_12_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_12_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_12_upstream_arb_share_counter_next_value);
  --cpu/instruction_master niosII_system_burst_12/upstream arbiterlock2, which is an e_assign
  cpu_instruction_master_arbiterlock2 <= niosII_system_burst_12_upstream_slavearbiterlockenable2 AND cpu_instruction_master_continuerequest;
  --niosII_system_burst_12_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_12_upstream_any_continuerequest <= std_logic'('1');
  --cpu_instruction_master_continuerequest continued request, which is an e_assign
  cpu_instruction_master_continuerequest <= std_logic'('1');
  internal_cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_12_upstream AND NOT ((cpu_instruction_master_read AND (((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_latency_counter))))))) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register)))));
  --unique name for niosII_system_burst_12_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_12_upstream_move_on_to_next_transaction <= niosII_system_burst_12_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_12_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_12_upstream, which is an e_mux
  niosII_system_burst_12_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_niosII_system_burst_12_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_instruction_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 6);
  --burstcount_fifo_for_niosII_system_burst_12_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_12_upstream : burstcount_fifo_for_niosII_system_burst_12_upstream_module
    port map(
      data_out => niosII_system_burst_12_upstream_transaction_burst_count,
      empty => niosII_system_burst_12_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input24,
      clk => clk,
      data_in => niosII_system_burst_12_upstream_selected_burstcount,
      read => niosII_system_burst_12_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input25,
      write => module_input26
    );

  module_input24 <= std_logic'('0');
  module_input25 <= std_logic'('0');
  module_input26 <= ((in_a_read_cycle AND NOT niosII_system_burst_12_upstream_waits_for_read) AND niosII_system_burst_12_upstream_load_fifo) AND NOT ((niosII_system_burst_12_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_12_upstream_burstcount_fifo_empty));

  --niosII_system_burst_12_upstream current burst minus one, which is an e_assign
  niosII_system_burst_12_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_12_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 6);
  --what to load in current_burst, for niosII_system_burst_12_upstream, which is an e_mux
  niosII_system_burst_12_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_12_upstream_waits_for_read)) AND NOT niosII_system_burst_12_upstream_load_fifo))) = '1'), (niosII_system_burst_12_upstream_selected_burstcount & std_logic_vector'("00")), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_12_upstream_waits_for_read) AND niosII_system_burst_12_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_12_upstream_burstcount_fifo_empty))) = '1'), (niosII_system_burst_12_upstream_selected_burstcount & std_logic_vector'("00")), A_WE_StdLogicVector((std_logic'((niosII_system_burst_12_upstream_this_cycle_is_the_last_burst)) = '1'), (niosII_system_burst_12_upstream_transaction_burst_count & std_logic_vector'("00")), (std_logic_vector'("00") & (niosII_system_burst_12_upstream_current_burst_minus_one))))), 6);
  --the current burst count for niosII_system_burst_12_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_12_upstream_current_burst <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_12_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_12_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_12_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_12_upstream_current_burst <= niosII_system_burst_12_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_12_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_12_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_12_upstream_waits_for_read)) AND niosII_system_burst_12_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_12_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_12_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_12_upstream_waits_for_read)) AND NOT niosII_system_burst_12_upstream_load_fifo) OR niosII_system_burst_12_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_12_upstream_load_fifo <= p0_niosII_system_burst_12_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_12_upstream, which is an e_assign
  niosII_system_burst_12_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_12_upstream_current_burst_minus_one)) AND niosII_system_burst_12_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_12_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_12_upstream : rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_12_upstream_module
    port map(
      data_out => cpu_instruction_master_rdv_fifo_output_from_niosII_system_burst_12_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_12_upstream,
      full => open,
      clear_fifo => module_input27,
      clk => clk,
      data_in => internal_cpu_instruction_master_granted_niosII_system_burst_12_upstream,
      read => niosII_system_burst_12_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input28,
      write => module_input29
    );

  module_input27 <= std_logic'('0');
  module_input28 <= std_logic'('0');
  module_input29 <= in_a_read_cycle AND NOT niosII_system_burst_12_upstream_waits_for_read;

  cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register <= NOT cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_12_upstream;
  --local readdatavalid cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream, which is an e_mux
  cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream <= niosII_system_burst_12_upstream_readdatavalid_from_sa;
  --byteaddress mux for niosII_system_burst_12/upstream, which is an e_mux
  niosII_system_burst_12_upstream_byteaddress <= cpu_instruction_master_address_to_slave (21 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_instruction_master_granted_niosII_system_burst_12_upstream <= internal_cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream;
  --cpu/instruction_master saved-grant niosII_system_burst_12/upstream, which is an e_assign
  cpu_instruction_master_saved_grant_niosII_system_burst_12_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_12_upstream;
  --allow new arb cycle for niosII_system_burst_12/upstream, which is an e_assign
  niosII_system_burst_12_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_12_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_12_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_12_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_12_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_12_upstream_begins_xfer) = '1'), niosII_system_burst_12_upstream_unreg_firsttransfer, niosII_system_burst_12_upstream_reg_firsttransfer);
  --niosII_system_burst_12_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_12_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_12_upstream_slavearbiterlockenable AND niosII_system_burst_12_upstream_any_continuerequest));
  --niosII_system_burst_12_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_12_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_12_upstream_begins_xfer) = '1' then 
        niosII_system_burst_12_upstream_reg_firsttransfer <= niosII_system_burst_12_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_12_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_12_upstream_beginbursttransfer_internal <= niosII_system_burst_12_upstream_begins_xfer;
  --niosII_system_burst_12_upstream_read assignment, which is an e_mux
  niosII_system_burst_12_upstream_read <= internal_cpu_instruction_master_granted_niosII_system_burst_12_upstream AND cpu_instruction_master_read;
  --niosII_system_burst_12_upstream_write assignment, which is an e_mux
  niosII_system_burst_12_upstream_write <= std_logic'('0');
  --niosII_system_burst_12_upstream_address mux, which is an e_mux
  niosII_system_burst_12_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & cpu_instruction_master_dbs_address(1 DOWNTO 0)), 22);
  --d1_niosII_system_burst_12_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_12_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_12_upstream_end_xfer <= niosII_system_burst_12_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_12_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_12_upstream_waits_for_read <= niosII_system_burst_12_upstream_in_a_read_cycle AND internal_niosII_system_burst_12_upstream_waitrequest_from_sa;
  --niosII_system_burst_12_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_12_upstream_in_a_read_cycle <= internal_cpu_instruction_master_granted_niosII_system_burst_12_upstream AND cpu_instruction_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_12_upstream_in_a_read_cycle;
  --niosII_system_burst_12_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_12_upstream_waits_for_write <= niosII_system_burst_12_upstream_in_a_write_cycle AND internal_niosII_system_burst_12_upstream_waitrequest_from_sa;
  --niosII_system_burst_12_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_12_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_12_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_12_upstream_counter <= std_logic'('0');
  --niosII_system_burst_12_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_12_upstream_byteenable <= Vector_To_Std_Logic(-SIGNED(std_logic_vector'("00000000000000000000000000000001")));
  --debugaccess mux, which is an e_mux
  niosII_system_burst_12_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_instruction_master_granted_niosII_system_burst_12_upstream <= internal_cpu_instruction_master_granted_niosII_system_burst_12_upstream;
  --vhdl renameroo for output signals
  cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream <= internal_cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream;
  --vhdl renameroo for output signals
  cpu_instruction_master_requests_niosII_system_burst_12_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_12_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_12_upstream_waitrequest_from_sa <= internal_niosII_system_burst_12_upstream_waitrequest_from_sa;
--synthesis translate_off
    --niosII_system_burst_12/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/instruction_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line59 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_instruction_master_requests_niosII_system_burst_12_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_instruction_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line59, now);
          write(write_line59, string'(": "));
          write(write_line59, string'("cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_12/upstream"));
          write(output, write_line59.all);
          deallocate (write_line59);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_12_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_tri_state_bridge_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal ext_flash_s1_wait_counter_eq_0 : IN STD_LOGIC;
                 signal incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_12_downstream_address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal niosII_system_burst_12_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_byteenable : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_granted_ext_flash_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_requests_ext_flash_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_12_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal niosII_system_burst_12_downstream_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_12_downstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_12_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_12_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_12_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_12_downstream_arbitrator;


architecture europa of niosII_system_burst_12_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_12_downstream_address_to_slave :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal internal_niosII_system_burst_12_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_niosII_system_burst_12_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_12_downstream_address_last_time :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_12_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_byteenable_last_time :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_is_granted_some_slave :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_niosII_system_burst_12_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pre_flush_niosII_system_burst_12_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 OR NOT niosII_system_burst_12_downstream_requests_ext_flash_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_12_downstream_granted_ext_flash_s1 OR NOT niosII_system_burst_12_downstream_qualified_request_ext_flash_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 OR NOT niosII_system_burst_12_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ext_flash_s1_wait_counter_eq_0 AND NOT d1_tri_state_bridge_avalon_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_12_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 OR NOT niosII_system_burst_12_downstream_write)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ext_flash_s1_wait_counter_eq_0 AND NOT d1_tri_state_bridge_avalon_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_12_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_12_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_12_downstream_address_to_slave <= niosII_system_burst_12_downstream_address;
  --niosII_system_burst_12_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_12_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_12_downstream_read_but_no_slave_selected <= (niosII_system_burst_12_downstream_read AND niosII_system_burst_12_downstream_run) AND NOT niosII_system_burst_12_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  niosII_system_burst_12_downstream_is_granted_some_slave <= niosII_system_burst_12_downstream_granted_ext_flash_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_12_downstream_readdatavalid <= niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_12_downstream_readdatavalid <= niosII_system_burst_12_downstream_read_but_no_slave_selected OR pre_flush_niosII_system_burst_12_downstream_readdatavalid;
  --niosII_system_burst_12/downstream readdata mux, which is an e_mux
  niosII_system_burst_12_downstream_readdata <= incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_12_downstream_waitrequest <= NOT niosII_system_burst_12_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_niosII_system_burst_12_downstream_latency_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      internal_niosII_system_burst_12_downstream_latency_counter <= p1_niosII_system_burst_12_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_niosII_system_burst_12_downstream_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((niosII_system_burst_12_downstream_run AND niosII_system_burst_12_downstream_read))) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_niosII_system_burst_12_downstream_latency_counter)) /= std_logic_vector'("00")), ((std_logic_vector'("0000000000000000000000000000000") & (internal_niosII_system_burst_12_downstream_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (A_REP(niosII_system_burst_12_downstream_requests_ext_flash_s1, 2))) AND std_logic_vector'("00000000000000000000000000000010")), 2);
  --niosII_system_burst_12_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_12_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_12_downstream_address_to_slave <= internal_niosII_system_burst_12_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_12_downstream_latency_counter <= internal_niosII_system_burst_12_downstream_latency_counter;
  --vhdl renameroo for output signals
  niosII_system_burst_12_downstream_waitrequest <= internal_niosII_system_burst_12_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_12_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_12_downstream_address_last_time <= std_logic_vector'("0000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_12_downstream_address_last_time <= niosII_system_burst_12_downstream_address;
      end if;

    end process;

    --niosII_system_burst_12/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_12_downstream_waitrequest AND ((niosII_system_burst_12_downstream_read OR niosII_system_burst_12_downstream_write));
      end if;

    end process;

    --niosII_system_burst_12_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line60 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_12_downstream_address /= niosII_system_burst_12_downstream_address_last_time))))) = '1' then 
          write(write_line60, now);
          write(write_line60, string'(": "));
          write(write_line60, string'("niosII_system_burst_12_downstream_address did not heed wait!!!"));
          write(output, write_line60.all);
          deallocate (write_line60);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_12_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_12_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_12_downstream_burstcount_last_time <= niosII_system_burst_12_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_12_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line61 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_12_downstream_burstcount) /= std_logic'(niosII_system_burst_12_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line61, now);
          write(write_line61, string'(": "));
          write(write_line61, string'("niosII_system_burst_12_downstream_burstcount did not heed wait!!!"));
          write(output, write_line61.all);
          deallocate (write_line61);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_12_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_12_downstream_byteenable_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_12_downstream_byteenable_last_time <= niosII_system_burst_12_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_12_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line62 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_12_downstream_byteenable) /= std_logic'(niosII_system_burst_12_downstream_byteenable_last_time)))))) = '1' then 
          write(write_line62, now);
          write(write_line62, string'(": "));
          write(write_line62, string'("niosII_system_burst_12_downstream_byteenable did not heed wait!!!"));
          write(output, write_line62.all);
          deallocate (write_line62);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_12_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_12_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_12_downstream_read_last_time <= niosII_system_burst_12_downstream_read;
      end if;

    end process;

    --niosII_system_burst_12_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line63 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_12_downstream_read) /= std_logic'(niosII_system_burst_12_downstream_read_last_time)))))) = '1' then 
          write(write_line63, now);
          write(write_line63, string'(": "));
          write(write_line63, string'("niosII_system_burst_12_downstream_read did not heed wait!!!"));
          write(output, write_line63.all);
          deallocate (write_line63);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_12_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_12_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_12_downstream_write_last_time <= niosII_system_burst_12_downstream_write;
      end if;

    end process;

    --niosII_system_burst_12_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line64 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_12_downstream_write) /= std_logic'(niosII_system_burst_12_downstream_write_last_time)))))) = '1' then 
          write(write_line64, now);
          write(write_line64, string'(": "));
          write(write_line64, string'("niosII_system_burst_12_downstream_write did not heed wait!!!"));
          write(output, write_line64.all);
          deallocate (write_line64);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_12_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_12_downstream_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_12_downstream_writedata_last_time <= niosII_system_burst_12_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_12_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line65 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_12_downstream_writedata /= niosII_system_burst_12_downstream_writedata_last_time)))) AND niosII_system_burst_12_downstream_write)) = '1' then 
          write(write_line65, now);
          write(write_line65, string'(": "));
          write(write_line65, string'("niosII_system_burst_12_downstream_writedata did not heed wait!!!"));
          write(output, write_line65.all);
          deallocate (write_line65);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_13_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_13_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_13_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("000000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("000000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("000000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("000000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_13_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_13_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_13_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_13_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal niosII_system_burst_13_upstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_13_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_13_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_byteenable_niosII_system_burst_13_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_granted_niosII_system_burst_13_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_13_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_13_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_13_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_13_upstream_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal niosII_system_burst_13_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_13_upstream_byteaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal niosII_system_burst_13_upstream_byteenable : OUT STD_LOGIC;
                 signal niosII_system_burst_13_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_13_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_13_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_13_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_13_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_13_upstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity niosII_system_burst_13_upstream_arbitrator;


architecture europa of niosII_system_burst_13_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_13_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_13_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_13_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_13_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_0 :  STD_LOGIC;
                signal cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_1 :  STD_LOGIC;
                signal cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_2 :  STD_LOGIC;
                signal cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_3 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_byteenable_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_13_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_13_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_13_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_13_upstream_write :  STD_LOGIC;
                signal module_input30 :  STD_LOGIC;
                signal module_input31 :  STD_LOGIC;
                signal module_input32 :  STD_LOGIC;
                signal module_input33 :  STD_LOGIC;
                signal module_input34 :  STD_LOGIC;
                signal module_input35 :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_13_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_13_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_13_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_13_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_current_burst :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_13_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_13_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_13_upstream_next_burst_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_13_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_selected_burstcount :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_13_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_13_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_13_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_13_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_13_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_13_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_13_upstream);
  --assign niosII_system_burst_13_upstream_readdatavalid_from_sa = niosII_system_burst_13_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_13_upstream_readdatavalid_from_sa <= niosII_system_burst_13_upstream_readdatavalid;
  --assign niosII_system_burst_13_upstream_readdata_from_sa = niosII_system_burst_13_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_13_upstream_readdata_from_sa <= niosII_system_burst_13_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_13_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 22) & std_logic_vector'("0000000000000000000000")) = std_logic_vector'("1010000000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_13_upstream_waitrequest_from_sa = niosII_system_burst_13_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_13_upstream_waitrequest_from_sa <= niosII_system_burst_13_upstream_waitrequest;
  --niosII_system_burst_13_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_13_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_13_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (A_SLL(cpu_data_master_burstcount,std_logic_vector'("00000000000000000000000000000010")))), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_13_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_13_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_13_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_13_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_13_upstream;
  --niosII_system_burst_13_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_13_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_13_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_13_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_13_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_13_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_13_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_13_upstream_allgrants <= niosII_system_burst_13_upstream_grant_vector;
  --niosII_system_burst_13_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_13_upstream_end_xfer <= NOT ((niosII_system_burst_13_upstream_waits_for_read OR niosII_system_burst_13_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_13_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_13_upstream <= niosII_system_burst_13_upstream_end_xfer AND (((NOT niosII_system_burst_13_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_13_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_13_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_13_upstream AND niosII_system_burst_13_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_13_upstream AND NOT niosII_system_burst_13_upstream_non_bursting_master_requests));
  --niosII_system_burst_13_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_13_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_13_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_13_upstream_arb_share_counter <= niosII_system_burst_13_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_13_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_13_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_13_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_13_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_13_upstream AND NOT niosII_system_burst_13_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_13_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_13_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_13/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_13_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_13_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_13_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_13_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_13/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_13_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_13_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_13_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_13_upstream <= internal_cpu_data_master_requests_niosII_system_burst_13_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_13_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_13_upstream_move_on_to_next_transaction <= niosII_system_burst_13_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_13_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_13_upstream, which is an e_mux
  niosII_system_burst_13_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_13_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 6);
  --burstcount_fifo_for_niosII_system_burst_13_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_13_upstream : burstcount_fifo_for_niosII_system_burst_13_upstream_module
    port map(
      data_out => niosII_system_burst_13_upstream_transaction_burst_count,
      empty => niosII_system_burst_13_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input30,
      clk => clk,
      data_in => niosII_system_burst_13_upstream_selected_burstcount,
      read => niosII_system_burst_13_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input31,
      write => module_input32
    );

  module_input30 <= std_logic'('0');
  module_input31 <= std_logic'('0');
  module_input32 <= ((in_a_read_cycle AND NOT niosII_system_burst_13_upstream_waits_for_read) AND niosII_system_burst_13_upstream_load_fifo) AND NOT ((niosII_system_burst_13_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_13_upstream_burstcount_fifo_empty));

  --niosII_system_burst_13_upstream current burst minus one, which is an e_assign
  niosII_system_burst_13_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_13_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 6);
  --what to load in current_burst, for niosII_system_burst_13_upstream, which is an e_mux
  niosII_system_burst_13_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_13_upstream_waits_for_read)) AND NOT niosII_system_burst_13_upstream_load_fifo))) = '1'), (niosII_system_burst_13_upstream_selected_burstcount & std_logic_vector'("00")), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_13_upstream_waits_for_read) AND niosII_system_burst_13_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_13_upstream_burstcount_fifo_empty))) = '1'), (niosII_system_burst_13_upstream_selected_burstcount & std_logic_vector'("00")), A_WE_StdLogicVector((std_logic'((niosII_system_burst_13_upstream_this_cycle_is_the_last_burst)) = '1'), (niosII_system_burst_13_upstream_transaction_burst_count & std_logic_vector'("00")), (std_logic_vector'("00") & (niosII_system_burst_13_upstream_current_burst_minus_one))))), 6);
  --the current burst count for niosII_system_burst_13_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_13_upstream_current_burst <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_13_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_13_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_13_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_13_upstream_current_burst <= niosII_system_burst_13_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_13_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_13_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_13_upstream_waits_for_read)) AND niosII_system_burst_13_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_13_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_13_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_13_upstream_waits_for_read)) AND NOT niosII_system_burst_13_upstream_load_fifo) OR niosII_system_burst_13_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_13_upstream_load_fifo <= p0_niosII_system_burst_13_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_13_upstream, which is an e_assign
  niosII_system_burst_13_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_13_upstream_current_burst_minus_one)) AND niosII_system_burst_13_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_13_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_13_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_13_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_13_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_13_upstream,
      full => open,
      clear_fifo => module_input33,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_13_upstream,
      read => niosII_system_burst_13_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input34,
      write => module_input35
    );

  module_input33 <= std_logic'('0');
  module_input34 <= std_logic'('0');
  module_input35 <= in_a_read_cycle AND NOT niosII_system_burst_13_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_13_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_13_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_13_upstream <= niosII_system_burst_13_upstream_readdatavalid_from_sa;
  --niosII_system_burst_13_upstream_writedata mux, which is an e_mux
  niosII_system_burst_13_upstream_writedata <= cpu_data_master_dbs_write_8;
  --byteaddress mux for niosII_system_burst_13/upstream, which is an e_mux
  niosII_system_burst_13_upstream_byteaddress <= cpu_data_master_address_to_slave (21 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_13_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_13_upstream;
  --cpu/data_master saved-grant niosII_system_burst_13/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_13_upstream <= internal_cpu_data_master_requests_niosII_system_burst_13_upstream;
  --allow new arb cycle for niosII_system_burst_13/upstream, which is an e_assign
  niosII_system_burst_13_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_13_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_13_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_13_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_13_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_13_upstream_begins_xfer) = '1'), niosII_system_burst_13_upstream_unreg_firsttransfer, niosII_system_burst_13_upstream_reg_firsttransfer);
  --niosII_system_burst_13_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_13_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_13_upstream_slavearbiterlockenable AND niosII_system_burst_13_upstream_any_continuerequest));
  --niosII_system_burst_13_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_13_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_13_upstream_begins_xfer) = '1' then 
        niosII_system_burst_13_upstream_reg_firsttransfer <= niosII_system_burst_13_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_13_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_13_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_13_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_13_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_13_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_13_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_13_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_13_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_13_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_13_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_13_upstream_begins_xfer) = '1' then 
        niosII_system_burst_13_upstream_bbt_burstcounter <= niosII_system_burst_13_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_13_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_13_upstream_beginbursttransfer_internal <= niosII_system_burst_13_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_13_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_13_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_13_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_13_upstream AND cpu_data_master_read;
  --niosII_system_burst_13_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_13_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_13_upstream AND cpu_data_master_write;
  --niosII_system_burst_13_upstream_address mux, which is an e_mux
  niosII_system_burst_13_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & cpu_data_master_dbs_address(1 DOWNTO 0)), 22);
  --d1_niosII_system_burst_13_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_13_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_13_upstream_end_xfer <= niosII_system_burst_13_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_13_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_13_upstream_waits_for_read <= niosII_system_burst_13_upstream_in_a_read_cycle AND internal_niosII_system_burst_13_upstream_waitrequest_from_sa;
  --niosII_system_burst_13_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_13_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_13_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_13_upstream_in_a_read_cycle;
  --niosII_system_burst_13_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_13_upstream_waits_for_write <= niosII_system_burst_13_upstream_in_a_write_cycle AND internal_niosII_system_burst_13_upstream_waitrequest_from_sa;
  --niosII_system_burst_13_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_13_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_13_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_13_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_13_upstream_counter <= std_logic'('0');
  --niosII_system_burst_13_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_13_upstream_byteenable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_13_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_cpu_data_master_byteenable_niosII_system_burst_13_upstream))), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  (cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_3, cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_2, cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_1, cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_0) <= cpu_data_master_byteenable;
  internal_cpu_data_master_byteenable_niosII_system_burst_13_upstream <= A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_0, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_1, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_2, cpu_data_master_byteenable_niosII_system_burst_13_upstream_segment_3)));
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_13_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_13_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_13_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_13_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_byteenable_niosII_system_burst_13_upstream <= internal_cpu_data_master_byteenable_niosII_system_burst_13_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_13_upstream <= internal_cpu_data_master_granted_niosII_system_burst_13_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_13_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_13_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_13_upstream <= internal_cpu_data_master_requests_niosII_system_burst_13_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_13_upstream_burstcount <= internal_niosII_system_burst_13_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_13_upstream_read <= internal_niosII_system_burst_13_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_13_upstream_waitrequest_from_sa <= internal_niosII_system_burst_13_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_13_upstream_write <= internal_niosII_system_burst_13_upstream_write;
--synthesis translate_off
    --niosII_system_burst_13/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line66 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_13_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line66, now);
          write(write_line66, string'(": "));
          write(write_line66, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_13/upstream"));
          write(output, write_line66.all);
          deallocate (write_line66);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_13_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_tri_state_bridge_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal ext_flash_s1_wait_counter_eq_0 : IN STD_LOGIC;
                 signal incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_13_downstream_address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal niosII_system_burst_13_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_byteenable : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_granted_ext_flash_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_requests_ext_flash_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_13_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal niosII_system_burst_13_downstream_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_13_downstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_13_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_13_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_13_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_13_downstream_arbitrator;


architecture europa of niosII_system_burst_13_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_13_downstream_address_to_slave :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal internal_niosII_system_burst_13_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_niosII_system_burst_13_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_13_downstream_address_last_time :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_13_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_byteenable_last_time :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_is_granted_some_slave :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_niosII_system_burst_13_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pre_flush_niosII_system_burst_13_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 OR NOT niosII_system_burst_13_downstream_requests_ext_flash_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_13_downstream_granted_ext_flash_s1 OR NOT niosII_system_burst_13_downstream_qualified_request_ext_flash_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 OR NOT niosII_system_burst_13_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ext_flash_s1_wait_counter_eq_0 AND NOT d1_tri_state_bridge_avalon_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_13_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 OR NOT niosII_system_burst_13_downstream_write)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ext_flash_s1_wait_counter_eq_0 AND NOT d1_tri_state_bridge_avalon_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_13_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_13_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_13_downstream_address_to_slave <= niosII_system_burst_13_downstream_address;
  --niosII_system_burst_13_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_13_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_13_downstream_read_but_no_slave_selected <= (niosII_system_burst_13_downstream_read AND niosII_system_burst_13_downstream_run) AND NOT niosII_system_burst_13_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  niosII_system_burst_13_downstream_is_granted_some_slave <= niosII_system_burst_13_downstream_granted_ext_flash_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_13_downstream_readdatavalid <= niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_13_downstream_readdatavalid <= niosII_system_burst_13_downstream_read_but_no_slave_selected OR pre_flush_niosII_system_burst_13_downstream_readdatavalid;
  --niosII_system_burst_13/downstream readdata mux, which is an e_mux
  niosII_system_burst_13_downstream_readdata <= incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_13_downstream_waitrequest <= NOT niosII_system_burst_13_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_niosII_system_burst_13_downstream_latency_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      internal_niosII_system_burst_13_downstream_latency_counter <= p1_niosII_system_burst_13_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_niosII_system_burst_13_downstream_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((niosII_system_burst_13_downstream_run AND niosII_system_burst_13_downstream_read))) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_niosII_system_burst_13_downstream_latency_counter)) /= std_logic_vector'("00")), ((std_logic_vector'("0000000000000000000000000000000") & (internal_niosII_system_burst_13_downstream_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (A_REP(niosII_system_burst_13_downstream_requests_ext_flash_s1, 2))) AND std_logic_vector'("00000000000000000000000000000010")), 2);
  --niosII_system_burst_13_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_13_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_13_downstream_address_to_slave <= internal_niosII_system_burst_13_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_13_downstream_latency_counter <= internal_niosII_system_burst_13_downstream_latency_counter;
  --vhdl renameroo for output signals
  niosII_system_burst_13_downstream_waitrequest <= internal_niosII_system_burst_13_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_13_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_13_downstream_address_last_time <= std_logic_vector'("0000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_13_downstream_address_last_time <= niosII_system_burst_13_downstream_address;
      end if;

    end process;

    --niosII_system_burst_13/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_13_downstream_waitrequest AND ((niosII_system_burst_13_downstream_read OR niosII_system_burst_13_downstream_write));
      end if;

    end process;

    --niosII_system_burst_13_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line67 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_13_downstream_address /= niosII_system_burst_13_downstream_address_last_time))))) = '1' then 
          write(write_line67, now);
          write(write_line67, string'(": "));
          write(write_line67, string'("niosII_system_burst_13_downstream_address did not heed wait!!!"));
          write(output, write_line67.all);
          deallocate (write_line67);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_13_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_13_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_13_downstream_burstcount_last_time <= niosII_system_burst_13_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_13_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line68 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_13_downstream_burstcount) /= std_logic'(niosII_system_burst_13_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line68, now);
          write(write_line68, string'(": "));
          write(write_line68, string'("niosII_system_burst_13_downstream_burstcount did not heed wait!!!"));
          write(output, write_line68.all);
          deallocate (write_line68);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_13_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_13_downstream_byteenable_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_13_downstream_byteenable_last_time <= niosII_system_burst_13_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_13_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line69 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_13_downstream_byteenable) /= std_logic'(niosII_system_burst_13_downstream_byteenable_last_time)))))) = '1' then 
          write(write_line69, now);
          write(write_line69, string'(": "));
          write(write_line69, string'("niosII_system_burst_13_downstream_byteenable did not heed wait!!!"));
          write(output, write_line69.all);
          deallocate (write_line69);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_13_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_13_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_13_downstream_read_last_time <= niosII_system_burst_13_downstream_read;
      end if;

    end process;

    --niosII_system_burst_13_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line70 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_13_downstream_read) /= std_logic'(niosII_system_burst_13_downstream_read_last_time)))))) = '1' then 
          write(write_line70, now);
          write(write_line70, string'(": "));
          write(write_line70, string'("niosII_system_burst_13_downstream_read did not heed wait!!!"));
          write(output, write_line70.all);
          deallocate (write_line70);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_13_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_13_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_13_downstream_write_last_time <= niosII_system_burst_13_downstream_write;
      end if;

    end process;

    --niosII_system_burst_13_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line71 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_13_downstream_write) /= std_logic'(niosII_system_burst_13_downstream_write_last_time)))))) = '1' then 
          write(write_line71, now);
          write(write_line71, string'(": "));
          write(write_line71, string'("niosII_system_burst_13_downstream_write did not heed wait!!!"));
          write(output, write_line71.all);
          deallocate (write_line71);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_13_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_13_downstream_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_13_downstream_writedata_last_time <= niosII_system_burst_13_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_13_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line72 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_13_downstream_writedata /= niosII_system_burst_13_downstream_writedata_last_time)))) AND niosII_system_burst_13_downstream_write)) = '1' then 
          write(write_line72, now);
          write(write_line72, string'(": "));
          write(write_line72, string'("niosII_system_burst_13_downstream_writedata did not heed wait!!!"));
          write(output, write_line72.all);
          deallocate (write_line72);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_14_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_14_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_14_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_14_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_14_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_14_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_14_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_14_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_14_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_14_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_14_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_14_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_14_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_14_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_14_upstream_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_14_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_14_upstream_byteaddress : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_14_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_14_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_14_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_14_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_14_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_14_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_14_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity niosII_system_burst_14_upstream_arbitrator;


architecture europa of niosII_system_burst_14_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_14_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_14_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_14_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_14_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_14_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_14_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_14_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_14_upstream_write :  STD_LOGIC;
                signal module_input36 :  STD_LOGIC;
                signal module_input37 :  STD_LOGIC;
                signal module_input38 :  STD_LOGIC;
                signal module_input39 :  STD_LOGIC;
                signal module_input40 :  STD_LOGIC;
                signal module_input41 :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_14_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_14_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_14_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_14_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_14_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_14_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_14_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_14_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_14_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_14_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_14_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_14_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_14_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_14_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_14_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_14_upstream);
  --assign niosII_system_burst_14_upstream_readdatavalid_from_sa = niosII_system_burst_14_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_14_upstream_readdatavalid_from_sa <= niosII_system_burst_14_upstream_readdatavalid;
  --assign niosII_system_burst_14_upstream_readdata_from_sa = niosII_system_burst_14_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_14_upstream_readdata_from_sa <= niosII_system_burst_14_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_14_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1100100001001000011000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_14_upstream_waitrequest_from_sa = niosII_system_burst_14_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_14_upstream_waitrequest_from_sa <= niosII_system_burst_14_upstream_waitrequest;
  --niosII_system_burst_14_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_14_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_14_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_14_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_14_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_14_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_14_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_14_upstream;
  --niosII_system_burst_14_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_14_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_14_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_14_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_14_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_14_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_14_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_14_upstream_allgrants <= niosII_system_burst_14_upstream_grant_vector;
  --niosII_system_burst_14_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_14_upstream_end_xfer <= NOT ((niosII_system_burst_14_upstream_waits_for_read OR niosII_system_burst_14_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_14_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_14_upstream <= niosII_system_burst_14_upstream_end_xfer AND (((NOT niosII_system_burst_14_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_14_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_14_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_14_upstream AND niosII_system_burst_14_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_14_upstream AND NOT niosII_system_burst_14_upstream_non_bursting_master_requests));
  --niosII_system_burst_14_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_14_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_14_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_14_upstream_arb_share_counter <= niosII_system_burst_14_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_14_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_14_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_14_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_14_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_14_upstream AND NOT niosII_system_burst_14_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_14_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_14_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_14/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_14_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_14_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_14_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_14_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_14/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_14_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_14_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_14_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_14_upstream <= internal_cpu_data_master_requests_niosII_system_burst_14_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_14_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_14_upstream_move_on_to_next_transaction <= niosII_system_burst_14_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_14_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_14_upstream, which is an e_mux
  niosII_system_burst_14_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_14_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_14_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_14_upstream : burstcount_fifo_for_niosII_system_burst_14_upstream_module
    port map(
      data_out => niosII_system_burst_14_upstream_transaction_burst_count,
      empty => niosII_system_burst_14_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input36,
      clk => clk,
      data_in => niosII_system_burst_14_upstream_selected_burstcount,
      read => niosII_system_burst_14_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input37,
      write => module_input38
    );

  module_input36 <= std_logic'('0');
  module_input37 <= std_logic'('0');
  module_input38 <= ((in_a_read_cycle AND NOT niosII_system_burst_14_upstream_waits_for_read) AND niosII_system_burst_14_upstream_load_fifo) AND NOT ((niosII_system_burst_14_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_14_upstream_burstcount_fifo_empty));

  --niosII_system_burst_14_upstream current burst minus one, which is an e_assign
  niosII_system_burst_14_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_14_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_14_upstream, which is an e_mux
  niosII_system_burst_14_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_14_upstream_waits_for_read)) AND NOT niosII_system_burst_14_upstream_load_fifo))) = '1'), niosII_system_burst_14_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_14_upstream_waits_for_read) AND niosII_system_burst_14_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_14_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_14_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_14_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_14_upstream_transaction_burst_count, niosII_system_burst_14_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_14_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_14_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_14_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_14_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_14_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_14_upstream_current_burst <= niosII_system_burst_14_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_14_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_14_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_14_upstream_waits_for_read)) AND niosII_system_burst_14_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_14_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_14_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_14_upstream_waits_for_read)) AND NOT niosII_system_burst_14_upstream_load_fifo) OR niosII_system_burst_14_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_14_upstream_load_fifo <= p0_niosII_system_burst_14_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_14_upstream, which is an e_assign
  niosII_system_burst_14_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_14_upstream_current_burst_minus_one)) AND niosII_system_burst_14_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_14_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_14_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_14_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_14_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_14_upstream,
      full => open,
      clear_fifo => module_input39,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_14_upstream,
      read => niosII_system_burst_14_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input40,
      write => module_input41
    );

  module_input39 <= std_logic'('0');
  module_input40 <= std_logic'('0');
  module_input41 <= in_a_read_cycle AND NOT niosII_system_burst_14_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_14_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_14_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_14_upstream <= niosII_system_burst_14_upstream_readdatavalid_from_sa;
  --niosII_system_burst_14_upstream_writedata mux, which is an e_mux
  niosII_system_burst_14_upstream_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --byteaddress mux for niosII_system_burst_14/upstream, which is an e_mux
  niosII_system_burst_14_upstream_byteaddress <= cpu_data_master_address_to_slave (3 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_14_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_14_upstream;
  --cpu/data_master saved-grant niosII_system_burst_14/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_14_upstream <= internal_cpu_data_master_requests_niosII_system_burst_14_upstream;
  --allow new arb cycle for niosII_system_burst_14/upstream, which is an e_assign
  niosII_system_burst_14_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_14_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_14_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_14_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_14_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_14_upstream_begins_xfer) = '1'), niosII_system_burst_14_upstream_unreg_firsttransfer, niosII_system_burst_14_upstream_reg_firsttransfer);
  --niosII_system_burst_14_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_14_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_14_upstream_slavearbiterlockenable AND niosII_system_burst_14_upstream_any_continuerequest));
  --niosII_system_burst_14_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_14_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_14_upstream_begins_xfer) = '1' then 
        niosII_system_burst_14_upstream_reg_firsttransfer <= niosII_system_burst_14_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_14_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_14_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_14_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_14_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_14_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_14_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_14_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_14_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_14_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_14_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_14_upstream_begins_xfer) = '1' then 
        niosII_system_burst_14_upstream_bbt_burstcounter <= niosII_system_burst_14_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_14_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_14_upstream_beginbursttransfer_internal <= niosII_system_burst_14_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_14_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_14_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_14_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_14_upstream AND cpu_data_master_read;
  --niosII_system_burst_14_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_14_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_14_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_14_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_14_upstream_address mux, which is an e_mux
  niosII_system_burst_14_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_14_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_niosII_system_burst_14_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_14_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_14_upstream_end_xfer <= niosII_system_burst_14_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_14_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_14_upstream_waits_for_read <= niosII_system_burst_14_upstream_in_a_read_cycle AND internal_niosII_system_burst_14_upstream_waitrequest_from_sa;
  --niosII_system_burst_14_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_14_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_14_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_14_upstream_in_a_read_cycle;
  --niosII_system_burst_14_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_14_upstream_waits_for_write <= niosII_system_burst_14_upstream_in_a_write_cycle AND internal_niosII_system_burst_14_upstream_waitrequest_from_sa;
  --niosII_system_burst_14_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_14_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_14_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_14_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_14_upstream_counter <= std_logic'('0');
  --niosII_system_burst_14_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_14_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_14_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_14_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_14_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_14_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_14_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_14_upstream <= internal_cpu_data_master_granted_niosII_system_burst_14_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_14_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_14_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_14_upstream <= internal_cpu_data_master_requests_niosII_system_burst_14_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_14_upstream_burstcount <= internal_niosII_system_burst_14_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_14_upstream_read <= internal_niosII_system_burst_14_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_14_upstream_waitrequest_from_sa <= internal_niosII_system_burst_14_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_14_upstream_write <= internal_niosII_system_burst_14_upstream_write;
--synthesis translate_off
    --niosII_system_burst_14/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line73 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_14_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line73, now);
          write(write_line73, string'(": "));
          write(write_line73, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_14/upstream"));
          write(output, write_line73.all);
          deallocate (write_line73);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_14_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_seven_seg_pio_s1_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_14_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal seven_seg_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal niosII_system_burst_14_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_14_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_14_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_14_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_14_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_14_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_14_downstream_arbitrator;


architecture europa of niosII_system_burst_14_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_14_downstream_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_niosII_system_burst_14_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_address_last_time :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_14_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_14_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_flush_niosII_system_burst_14_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 OR NOT niosII_system_burst_14_downstream_requests_seven_seg_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 OR NOT niosII_system_burst_14_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_seven_seg_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_14_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 OR NOT niosII_system_burst_14_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_14_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_14_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_14_downstream_address_to_slave <= niosII_system_burst_14_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_14_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_14_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_14_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1)))));
  --niosII_system_burst_14/downstream readdata mux, which is an e_mux
  niosII_system_burst_14_downstream_readdata <= seven_seg_pio_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_14_downstream_waitrequest <= NOT niosII_system_burst_14_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_14_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_14_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_14_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_14_downstream_address_to_slave <= internal_niosII_system_burst_14_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_14_downstream_waitrequest <= internal_niosII_system_burst_14_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_14_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_14_downstream_address_last_time <= std_logic_vector'("000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_14_downstream_address_last_time <= niosII_system_burst_14_downstream_address;
      end if;

    end process;

    --niosII_system_burst_14/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_14_downstream_waitrequest AND ((niosII_system_burst_14_downstream_read OR niosII_system_burst_14_downstream_write));
      end if;

    end process;

    --niosII_system_burst_14_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line74 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_14_downstream_address /= niosII_system_burst_14_downstream_address_last_time))))) = '1' then 
          write(write_line74, now);
          write(write_line74, string'(": "));
          write(write_line74, string'("niosII_system_burst_14_downstream_address did not heed wait!!!"));
          write(output, write_line74.all);
          deallocate (write_line74);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_14_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_14_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_14_downstream_burstcount_last_time <= niosII_system_burst_14_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_14_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line75 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_14_downstream_burstcount) /= std_logic'(niosII_system_burst_14_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line75, now);
          write(write_line75, string'(": "));
          write(write_line75, string'("niosII_system_burst_14_downstream_burstcount did not heed wait!!!"));
          write(output, write_line75.all);
          deallocate (write_line75);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_14_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_14_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_14_downstream_byteenable_last_time <= niosII_system_burst_14_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_14_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line76 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_14_downstream_byteenable /= niosII_system_burst_14_downstream_byteenable_last_time))))) = '1' then 
          write(write_line76, now);
          write(write_line76, string'(": "));
          write(write_line76, string'("niosII_system_burst_14_downstream_byteenable did not heed wait!!!"));
          write(output, write_line76.all);
          deallocate (write_line76);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_14_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_14_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_14_downstream_read_last_time <= niosII_system_burst_14_downstream_read;
      end if;

    end process;

    --niosII_system_burst_14_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line77 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_14_downstream_read) /= std_logic'(niosII_system_burst_14_downstream_read_last_time)))))) = '1' then 
          write(write_line77, now);
          write(write_line77, string'(": "));
          write(write_line77, string'("niosII_system_burst_14_downstream_read did not heed wait!!!"));
          write(output, write_line77.all);
          deallocate (write_line77);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_14_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_14_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_14_downstream_write_last_time <= niosII_system_burst_14_downstream_write;
      end if;

    end process;

    --niosII_system_burst_14_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line78 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_14_downstream_write) /= std_logic'(niosII_system_burst_14_downstream_write_last_time)))))) = '1' then 
          write(write_line78, now);
          write(write_line78, string'(": "));
          write(write_line78, string'("niosII_system_burst_14_downstream_write did not heed wait!!!"));
          write(output, write_line78.all);
          deallocate (write_line78);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_14_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_14_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_14_downstream_writedata_last_time <= niosII_system_burst_14_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_14_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line79 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_14_downstream_writedata /= niosII_system_burst_14_downstream_writedata_last_time)))) AND niosII_system_burst_14_downstream_write)) = '1' then 
          write(write_line79, now);
          write(write_line79, string'(": "));
          write(write_line79, string'("niosII_system_burst_14_downstream_writedata did not heed wait!!!"));
          write(output, write_line79.all);
          deallocate (write_line79);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_15_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_15_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_15_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_15_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_15_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_15_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_15_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_15_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_15_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_15_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_15_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_15_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_15_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_15_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_15_upstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_15_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_15_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_15_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_15_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_15_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_15_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_15_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_15_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_15_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity niosII_system_burst_15_upstream_arbitrator;


architecture europa of niosII_system_burst_15_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_15_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_15_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_15_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_15_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_15_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_15_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_15_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_15_upstream_write :  STD_LOGIC;
                signal module_input42 :  STD_LOGIC;
                signal module_input43 :  STD_LOGIC;
                signal module_input44 :  STD_LOGIC;
                signal module_input45 :  STD_LOGIC;
                signal module_input46 :  STD_LOGIC;
                signal module_input47 :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_15_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_15_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_15_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_15_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_15_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_15_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_15_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_15_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_15_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_15_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_15_upstream);
  --assign niosII_system_burst_15_upstream_readdatavalid_from_sa = niosII_system_burst_15_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_15_upstream_readdatavalid_from_sa <= niosII_system_burst_15_upstream_readdatavalid;
  --assign niosII_system_burst_15_upstream_readdata_from_sa = niosII_system_burst_15_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_15_upstream_readdata_from_sa <= niosII_system_burst_15_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_15_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1100100001001000000100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_15_upstream_waitrequest_from_sa = niosII_system_burst_15_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_15_upstream_waitrequest_from_sa <= niosII_system_burst_15_upstream_waitrequest;
  --niosII_system_burst_15_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_15_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_15_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_15_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_15_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_15_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_15_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_15_upstream;
  --niosII_system_burst_15_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_15_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_15_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_15_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_15_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_15_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_15_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_15_upstream_allgrants <= niosII_system_burst_15_upstream_grant_vector;
  --niosII_system_burst_15_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_15_upstream_end_xfer <= NOT ((niosII_system_burst_15_upstream_waits_for_read OR niosII_system_burst_15_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_15_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_15_upstream <= niosII_system_burst_15_upstream_end_xfer AND (((NOT niosII_system_burst_15_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_15_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_15_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_15_upstream AND niosII_system_burst_15_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_15_upstream AND NOT niosII_system_burst_15_upstream_non_bursting_master_requests));
  --niosII_system_burst_15_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_15_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_15_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_15_upstream_arb_share_counter <= niosII_system_burst_15_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_15_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_15_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_15_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_15_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_15_upstream AND NOT niosII_system_burst_15_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_15_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_15_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_15/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_15_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_15_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_15_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_15_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_15/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_15_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_15_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_15_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_15_upstream <= internal_cpu_data_master_requests_niosII_system_burst_15_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_15_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_15_upstream_move_on_to_next_transaction <= niosII_system_burst_15_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_15_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_15_upstream, which is an e_mux
  niosII_system_burst_15_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_15_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_15_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_15_upstream : burstcount_fifo_for_niosII_system_burst_15_upstream_module
    port map(
      data_out => niosII_system_burst_15_upstream_transaction_burst_count,
      empty => niosII_system_burst_15_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input42,
      clk => clk,
      data_in => niosII_system_burst_15_upstream_selected_burstcount,
      read => niosII_system_burst_15_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input43,
      write => module_input44
    );

  module_input42 <= std_logic'('0');
  module_input43 <= std_logic'('0');
  module_input44 <= ((in_a_read_cycle AND NOT niosII_system_burst_15_upstream_waits_for_read) AND niosII_system_burst_15_upstream_load_fifo) AND NOT ((niosII_system_burst_15_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_15_upstream_burstcount_fifo_empty));

  --niosII_system_burst_15_upstream current burst minus one, which is an e_assign
  niosII_system_burst_15_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_15_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_15_upstream, which is an e_mux
  niosII_system_burst_15_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_15_upstream_waits_for_read)) AND NOT niosII_system_burst_15_upstream_load_fifo))) = '1'), niosII_system_burst_15_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_15_upstream_waits_for_read) AND niosII_system_burst_15_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_15_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_15_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_15_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_15_upstream_transaction_burst_count, niosII_system_burst_15_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_15_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_15_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_15_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_15_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_15_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_15_upstream_current_burst <= niosII_system_burst_15_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_15_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_15_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_15_upstream_waits_for_read)) AND niosII_system_burst_15_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_15_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_15_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_15_upstream_waits_for_read)) AND NOT niosII_system_burst_15_upstream_load_fifo) OR niosII_system_burst_15_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_15_upstream_load_fifo <= p0_niosII_system_burst_15_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_15_upstream, which is an e_assign
  niosII_system_burst_15_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_15_upstream_current_burst_minus_one)) AND niosII_system_burst_15_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_15_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_15_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_15_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_15_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_15_upstream,
      full => open,
      clear_fifo => module_input45,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_15_upstream,
      read => niosII_system_burst_15_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input46,
      write => module_input47
    );

  module_input45 <= std_logic'('0');
  module_input46 <= std_logic'('0');
  module_input47 <= in_a_read_cycle AND NOT niosII_system_burst_15_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_15_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_15_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_15_upstream <= niosII_system_burst_15_upstream_readdatavalid_from_sa;
  --niosII_system_burst_15_upstream_writedata mux, which is an e_mux
  niosII_system_burst_15_upstream_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --byteaddress mux for niosII_system_burst_15/upstream, which is an e_mux
  niosII_system_burst_15_upstream_byteaddress <= cpu_data_master_address_to_slave (4 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_15_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_15_upstream;
  --cpu/data_master saved-grant niosII_system_burst_15/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_15_upstream <= internal_cpu_data_master_requests_niosII_system_burst_15_upstream;
  --allow new arb cycle for niosII_system_burst_15/upstream, which is an e_assign
  niosII_system_burst_15_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_15_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_15_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_15_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_15_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_15_upstream_begins_xfer) = '1'), niosII_system_burst_15_upstream_unreg_firsttransfer, niosII_system_burst_15_upstream_reg_firsttransfer);
  --niosII_system_burst_15_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_15_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_15_upstream_slavearbiterlockenable AND niosII_system_burst_15_upstream_any_continuerequest));
  --niosII_system_burst_15_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_15_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_15_upstream_begins_xfer) = '1' then 
        niosII_system_burst_15_upstream_reg_firsttransfer <= niosII_system_burst_15_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_15_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_15_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_15_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_15_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_15_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_15_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_15_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_15_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_15_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_15_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_15_upstream_begins_xfer) = '1' then 
        niosII_system_burst_15_upstream_bbt_burstcounter <= niosII_system_burst_15_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_15_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_15_upstream_beginbursttransfer_internal <= niosII_system_burst_15_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_15_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_15_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_15_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_15_upstream AND cpu_data_master_read;
  --niosII_system_burst_15_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_15_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_15_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_15_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_15_upstream_address mux, which is an e_mux
  niosII_system_burst_15_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_15_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --d1_niosII_system_burst_15_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_15_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_15_upstream_end_xfer <= niosII_system_burst_15_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_15_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_15_upstream_waits_for_read <= niosII_system_burst_15_upstream_in_a_read_cycle AND internal_niosII_system_burst_15_upstream_waitrequest_from_sa;
  --niosII_system_burst_15_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_15_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_15_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_15_upstream_in_a_read_cycle;
  --niosII_system_burst_15_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_15_upstream_waits_for_write <= niosII_system_burst_15_upstream_in_a_write_cycle AND internal_niosII_system_burst_15_upstream_waitrequest_from_sa;
  --niosII_system_burst_15_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_15_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_15_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_15_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_15_upstream_counter <= std_logic'('0');
  --niosII_system_burst_15_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_15_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_15_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_15_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_15_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_15_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_15_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_15_upstream <= internal_cpu_data_master_granted_niosII_system_burst_15_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_15_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_15_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_15_upstream <= internal_cpu_data_master_requests_niosII_system_burst_15_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_15_upstream_burstcount <= internal_niosII_system_burst_15_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_15_upstream_read <= internal_niosII_system_burst_15_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_15_upstream_waitrequest_from_sa <= internal_niosII_system_burst_15_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_15_upstream_write <= internal_niosII_system_burst_15_upstream_write;
--synthesis translate_off
    --niosII_system_burst_15/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line80 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_15_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line80, now);
          write(write_line80, string'(": "));
          write(write_line80, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_15/upstream"));
          write(output, write_line80.all);
          deallocate (write_line80);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_15_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_high_res_timer_s1_end_xfer : IN STD_LOGIC;
                 signal high_res_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_15_downstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_15_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_15_downstream_granted_high_res_timer_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_requests_high_res_timer_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_15_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_15_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_15_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_15_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_15_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_15_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_15_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_15_downstream_arbitrator;


architecture europa of niosII_system_burst_15_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_15_downstream_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_15_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_15_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_flush_niosII_system_burst_15_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 OR NOT niosII_system_burst_15_downstream_requests_high_res_timer_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 OR NOT niosII_system_burst_15_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_high_res_timer_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_15_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 OR NOT niosII_system_burst_15_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_15_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_15_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_15_downstream_address_to_slave <= niosII_system_burst_15_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_15_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_15_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_15_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1)))));
  --niosII_system_burst_15/downstream readdata mux, which is an e_mux
  niosII_system_burst_15_downstream_readdata <= high_res_timer_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_15_downstream_waitrequest <= NOT niosII_system_burst_15_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_15_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_15_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_15_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_15_downstream_address_to_slave <= internal_niosII_system_burst_15_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_15_downstream_waitrequest <= internal_niosII_system_burst_15_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_15_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_15_downstream_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_15_downstream_address_last_time <= niosII_system_burst_15_downstream_address;
      end if;

    end process;

    --niosII_system_burst_15/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_15_downstream_waitrequest AND ((niosII_system_burst_15_downstream_read OR niosII_system_burst_15_downstream_write));
      end if;

    end process;

    --niosII_system_burst_15_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line81 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_15_downstream_address /= niosII_system_burst_15_downstream_address_last_time))))) = '1' then 
          write(write_line81, now);
          write(write_line81, string'(": "));
          write(write_line81, string'("niosII_system_burst_15_downstream_address did not heed wait!!!"));
          write(output, write_line81.all);
          deallocate (write_line81);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_15_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_15_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_15_downstream_burstcount_last_time <= niosII_system_burst_15_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_15_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line82 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_15_downstream_burstcount) /= std_logic'(niosII_system_burst_15_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line82, now);
          write(write_line82, string'(": "));
          write(write_line82, string'("niosII_system_burst_15_downstream_burstcount did not heed wait!!!"));
          write(output, write_line82.all);
          deallocate (write_line82);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_15_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_15_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_15_downstream_byteenable_last_time <= niosII_system_burst_15_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_15_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line83 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_15_downstream_byteenable /= niosII_system_burst_15_downstream_byteenable_last_time))))) = '1' then 
          write(write_line83, now);
          write(write_line83, string'(": "));
          write(write_line83, string'("niosII_system_burst_15_downstream_byteenable did not heed wait!!!"));
          write(output, write_line83.all);
          deallocate (write_line83);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_15_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_15_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_15_downstream_read_last_time <= niosII_system_burst_15_downstream_read;
      end if;

    end process;

    --niosII_system_burst_15_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line84 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_15_downstream_read) /= std_logic'(niosII_system_burst_15_downstream_read_last_time)))))) = '1' then 
          write(write_line84, now);
          write(write_line84, string'(": "));
          write(write_line84, string'("niosII_system_burst_15_downstream_read did not heed wait!!!"));
          write(output, write_line84.all);
          deallocate (write_line84);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_15_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_15_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_15_downstream_write_last_time <= niosII_system_burst_15_downstream_write;
      end if;

    end process;

    --niosII_system_burst_15_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line85 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_15_downstream_write) /= std_logic'(niosII_system_burst_15_downstream_write_last_time)))))) = '1' then 
          write(write_line85, now);
          write(write_line85, string'(": "));
          write(write_line85, string'("niosII_system_burst_15_downstream_write did not heed wait!!!"));
          write(output, write_line85.all);
          deallocate (write_line85);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_15_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_15_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_15_downstream_writedata_last_time <= niosII_system_burst_15_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_15_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line86 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_15_downstream_writedata /= niosII_system_burst_15_downstream_writedata_last_time)))) AND niosII_system_burst_15_downstream_write)) = '1' then 
          write(write_line86, now);
          write(write_line86, string'(": "));
          write(write_line86, string'("niosII_system_burst_15_downstream_writedata did not heed wait!!!"));
          write(output, write_line86.all);
          deallocate (write_line86);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_16_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_16_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_16_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_16_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_16_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_16_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_16_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_16_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_16_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_16_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_16_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_16_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_16_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_16_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_16_upstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_16_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_16_upstream_byteaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_16_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_16_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_16_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_16_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_16_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_16_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_16_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity niosII_system_burst_16_upstream_arbitrator;


architecture europa of niosII_system_burst_16_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_16_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_16_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_16_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_16_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_16_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_16_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_16_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_16_upstream_write :  STD_LOGIC;
                signal module_input48 :  STD_LOGIC;
                signal module_input49 :  STD_LOGIC;
                signal module_input50 :  STD_LOGIC;
                signal module_input51 :  STD_LOGIC;
                signal module_input52 :  STD_LOGIC;
                signal module_input53 :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_16_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_16_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_16_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_16_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_16_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_16_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_16_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_16_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_16_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_16_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_16_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_16_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_16_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_16_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_16_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_16_upstream);
  --assign niosII_system_burst_16_upstream_readdatavalid_from_sa = niosII_system_burst_16_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_16_upstream_readdatavalid_from_sa <= niosII_system_burst_16_upstream_readdatavalid;
  --assign niosII_system_burst_16_upstream_readdata_from_sa = niosII_system_burst_16_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_16_upstream_readdata_from_sa <= niosII_system_burst_16_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_16_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("1100100001001000011100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_16_upstream_waitrequest_from_sa = niosII_system_burst_16_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_16_upstream_waitrequest_from_sa <= niosII_system_burst_16_upstream_waitrequest;
  --niosII_system_burst_16_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_16_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_16_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_16_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_16_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_16_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_16_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_16_upstream;
  --niosII_system_burst_16_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_16_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_16_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_16_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_16_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_16_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_16_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_16_upstream_allgrants <= niosII_system_burst_16_upstream_grant_vector;
  --niosII_system_burst_16_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_16_upstream_end_xfer <= NOT ((niosII_system_burst_16_upstream_waits_for_read OR niosII_system_burst_16_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_16_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_16_upstream <= niosII_system_burst_16_upstream_end_xfer AND (((NOT niosII_system_burst_16_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_16_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_16_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_16_upstream AND niosII_system_burst_16_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_16_upstream AND NOT niosII_system_burst_16_upstream_non_bursting_master_requests));
  --niosII_system_burst_16_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_16_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_16_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_16_upstream_arb_share_counter <= niosII_system_burst_16_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_16_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_16_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_16_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_16_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_16_upstream AND NOT niosII_system_burst_16_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_16_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_16_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_16/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_16_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_16_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_16_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_16_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_16/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_16_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_16_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_16_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_16_upstream <= internal_cpu_data_master_requests_niosII_system_burst_16_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_16_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_16_upstream_move_on_to_next_transaction <= niosII_system_burst_16_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_16_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_16_upstream, which is an e_mux
  niosII_system_burst_16_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_16_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_16_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_16_upstream : burstcount_fifo_for_niosII_system_burst_16_upstream_module
    port map(
      data_out => niosII_system_burst_16_upstream_transaction_burst_count,
      empty => niosII_system_burst_16_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input48,
      clk => clk,
      data_in => niosII_system_burst_16_upstream_selected_burstcount,
      read => niosII_system_burst_16_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input49,
      write => module_input50
    );

  module_input48 <= std_logic'('0');
  module_input49 <= std_logic'('0');
  module_input50 <= ((in_a_read_cycle AND NOT niosII_system_burst_16_upstream_waits_for_read) AND niosII_system_burst_16_upstream_load_fifo) AND NOT ((niosII_system_burst_16_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_16_upstream_burstcount_fifo_empty));

  --niosII_system_burst_16_upstream current burst minus one, which is an e_assign
  niosII_system_burst_16_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_16_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_16_upstream, which is an e_mux
  niosII_system_burst_16_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_16_upstream_waits_for_read)) AND NOT niosII_system_burst_16_upstream_load_fifo))) = '1'), niosII_system_burst_16_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_16_upstream_waits_for_read) AND niosII_system_burst_16_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_16_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_16_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_16_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_16_upstream_transaction_burst_count, niosII_system_burst_16_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_16_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_16_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_16_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_16_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_16_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_16_upstream_current_burst <= niosII_system_burst_16_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_16_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_16_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_16_upstream_waits_for_read)) AND niosII_system_burst_16_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_16_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_16_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_16_upstream_waits_for_read)) AND NOT niosII_system_burst_16_upstream_load_fifo) OR niosII_system_burst_16_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_16_upstream_load_fifo <= p0_niosII_system_burst_16_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_16_upstream, which is an e_assign
  niosII_system_burst_16_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_16_upstream_current_burst_minus_one)) AND niosII_system_burst_16_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_16_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_16_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_16_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_16_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_16_upstream,
      full => open,
      clear_fifo => module_input51,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_16_upstream,
      read => niosII_system_burst_16_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input52,
      write => module_input53
    );

  module_input51 <= std_logic'('0');
  module_input52 <= std_logic'('0');
  module_input53 <= in_a_read_cycle AND NOT niosII_system_burst_16_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_16_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_16_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_16_upstream <= niosII_system_burst_16_upstream_readdatavalid_from_sa;
  --niosII_system_burst_16_upstream_writedata mux, which is an e_mux
  niosII_system_burst_16_upstream_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --byteaddress mux for niosII_system_burst_16/upstream, which is an e_mux
  niosII_system_burst_16_upstream_byteaddress <= cpu_data_master_address_to_slave (2 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_16_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_16_upstream;
  --cpu/data_master saved-grant niosII_system_burst_16/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_16_upstream <= internal_cpu_data_master_requests_niosII_system_burst_16_upstream;
  --allow new arb cycle for niosII_system_burst_16/upstream, which is an e_assign
  niosII_system_burst_16_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_16_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_16_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_16_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_16_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_16_upstream_begins_xfer) = '1'), niosII_system_burst_16_upstream_unreg_firsttransfer, niosII_system_burst_16_upstream_reg_firsttransfer);
  --niosII_system_burst_16_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_16_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_16_upstream_slavearbiterlockenable AND niosII_system_burst_16_upstream_any_continuerequest));
  --niosII_system_burst_16_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_16_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_16_upstream_begins_xfer) = '1' then 
        niosII_system_burst_16_upstream_reg_firsttransfer <= niosII_system_burst_16_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_16_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_16_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_16_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_16_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_16_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_16_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_16_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_16_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_16_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_16_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_16_upstream_begins_xfer) = '1' then 
        niosII_system_burst_16_upstream_bbt_burstcounter <= niosII_system_burst_16_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_16_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_16_upstream_beginbursttransfer_internal <= niosII_system_burst_16_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_16_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_16_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_16_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_16_upstream AND cpu_data_master_read;
  --niosII_system_burst_16_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_16_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_16_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_16_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_16_upstream_address mux, which is an e_mux
  niosII_system_burst_16_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_16_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_niosII_system_burst_16_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_16_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_16_upstream_end_xfer <= niosII_system_burst_16_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_16_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_16_upstream_waits_for_read <= niosII_system_burst_16_upstream_in_a_read_cycle AND internal_niosII_system_burst_16_upstream_waitrequest_from_sa;
  --niosII_system_burst_16_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_16_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_16_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_16_upstream_in_a_read_cycle;
  --niosII_system_burst_16_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_16_upstream_waits_for_write <= niosII_system_burst_16_upstream_in_a_write_cycle AND internal_niosII_system_burst_16_upstream_waitrequest_from_sa;
  --niosII_system_burst_16_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_16_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_16_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_16_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_16_upstream_counter <= std_logic'('0');
  --niosII_system_burst_16_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_16_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_16_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_16_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_16_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_16_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_16_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_16_upstream <= internal_cpu_data_master_granted_niosII_system_burst_16_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_16_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_16_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_16_upstream <= internal_cpu_data_master_requests_niosII_system_burst_16_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_16_upstream_burstcount <= internal_niosII_system_burst_16_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_16_upstream_read <= internal_niosII_system_burst_16_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_16_upstream_waitrequest_from_sa <= internal_niosII_system_burst_16_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_16_upstream_write <= internal_niosII_system_burst_16_upstream_write;
--synthesis translate_off
    --niosII_system_burst_16/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line87 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_16_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line87, now);
          write(write_line87, string'(": "));
          write(write_line87, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_16/upstream"));
          write(output, write_line87.all);
          deallocate (write_line87);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_16_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_dm9000a_inst_avalon_slave_0_end_xfer : IN STD_LOGIC;
                 signal dm9000a_inst_avalon_slave_0_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_16_downstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_16_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0 : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_16_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_16_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_16_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_16_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_16_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_16_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_16_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_16_downstream_arbitrator;


architecture europa of niosII_system_burst_16_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_16_downstream_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_niosII_system_burst_16_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_16_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_16_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_flush_niosII_system_burst_16_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 OR NOT niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 OR NOT niosII_system_burst_16_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_dm9000a_inst_avalon_slave_0_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_16_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 OR NOT niosII_system_burst_16_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_16_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_16_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_16_downstream_address_to_slave <= niosII_system_burst_16_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_16_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_16_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_16_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0)))));
  --niosII_system_burst_16/downstream readdata mux, which is an e_mux
  niosII_system_burst_16_downstream_readdata <= dm9000a_inst_avalon_slave_0_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_16_downstream_waitrequest <= NOT niosII_system_burst_16_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_16_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_16_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_16_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_16_downstream_address_to_slave <= internal_niosII_system_burst_16_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_16_downstream_waitrequest <= internal_niosII_system_burst_16_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_16_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_16_downstream_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_16_downstream_address_last_time <= niosII_system_burst_16_downstream_address;
      end if;

    end process;

    --niosII_system_burst_16/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_16_downstream_waitrequest AND ((niosII_system_burst_16_downstream_read OR niosII_system_burst_16_downstream_write));
      end if;

    end process;

    --niosII_system_burst_16_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line88 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_16_downstream_address /= niosII_system_burst_16_downstream_address_last_time))))) = '1' then 
          write(write_line88, now);
          write(write_line88, string'(": "));
          write(write_line88, string'("niosII_system_burst_16_downstream_address did not heed wait!!!"));
          write(output, write_line88.all);
          deallocate (write_line88);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_16_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_16_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_16_downstream_burstcount_last_time <= niosII_system_burst_16_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_16_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line89 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_16_downstream_burstcount) /= std_logic'(niosII_system_burst_16_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line89, now);
          write(write_line89, string'(": "));
          write(write_line89, string'("niosII_system_burst_16_downstream_burstcount did not heed wait!!!"));
          write(output, write_line89.all);
          deallocate (write_line89);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_16_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_16_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_16_downstream_byteenable_last_time <= niosII_system_burst_16_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_16_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line90 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_16_downstream_byteenable /= niosII_system_burst_16_downstream_byteenable_last_time))))) = '1' then 
          write(write_line90, now);
          write(write_line90, string'(": "));
          write(write_line90, string'("niosII_system_burst_16_downstream_byteenable did not heed wait!!!"));
          write(output, write_line90.all);
          deallocate (write_line90);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_16_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_16_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_16_downstream_read_last_time <= niosII_system_burst_16_downstream_read;
      end if;

    end process;

    --niosII_system_burst_16_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line91 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_16_downstream_read) /= std_logic'(niosII_system_burst_16_downstream_read_last_time)))))) = '1' then 
          write(write_line91, now);
          write(write_line91, string'(": "));
          write(write_line91, string'("niosII_system_burst_16_downstream_read did not heed wait!!!"));
          write(output, write_line91.all);
          deallocate (write_line91);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_16_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_16_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_16_downstream_write_last_time <= niosII_system_burst_16_downstream_write;
      end if;

    end process;

    --niosII_system_burst_16_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line92 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_16_downstream_write) /= std_logic'(niosII_system_burst_16_downstream_write_last_time)))))) = '1' then 
          write(write_line92, now);
          write(write_line92, string'(": "));
          write(write_line92, string'("niosII_system_burst_16_downstream_write did not heed wait!!!"));
          write(output, write_line92.all);
          deallocate (write_line92);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_16_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_16_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_16_downstream_writedata_last_time <= niosII_system_burst_16_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_16_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line93 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_16_downstream_writedata /= niosII_system_burst_16_downstream_writedata_last_time)))) AND niosII_system_burst_16_downstream_write)) = '1' then 
          write(write_line93, now);
          write(write_line93, string'(": "));
          write(write_line93, string'("niosII_system_burst_16_downstream_writedata did not heed wait!!!"));
          write(output, write_line93.all);
          deallocate (write_line93);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_17_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_17_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_17_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_17_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_17_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_17_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_17_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_17_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_17_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_17_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_17_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_17_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_17_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_17_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_17_upstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_17_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_17_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_17_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_17_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_17_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_17_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_17_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_17_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_17_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity niosII_system_burst_17_upstream_arbitrator;


architecture europa of niosII_system_burst_17_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_17_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_17_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_17_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_17_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_17_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_17_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_17_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_17_upstream_write :  STD_LOGIC;
                signal module_input54 :  STD_LOGIC;
                signal module_input55 :  STD_LOGIC;
                signal module_input56 :  STD_LOGIC;
                signal module_input57 :  STD_LOGIC;
                signal module_input58 :  STD_LOGIC;
                signal module_input59 :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_17_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_17_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_17_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_17_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_17_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_17_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_17_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_17_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_17_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_17_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_17_upstream);
  --assign niosII_system_burst_17_upstream_readdatavalid_from_sa = niosII_system_burst_17_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_17_upstream_readdatavalid_from_sa <= niosII_system_burst_17_upstream_readdatavalid;
  --assign niosII_system_burst_17_upstream_readdata_from_sa = niosII_system_burst_17_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_17_upstream_readdata_from_sa <= niosII_system_burst_17_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_17_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1100100001001000001000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_17_upstream_waitrequest_from_sa = niosII_system_burst_17_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_17_upstream_waitrequest_from_sa <= niosII_system_burst_17_upstream_waitrequest;
  --niosII_system_burst_17_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_17_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_17_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_17_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_17_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_17_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_17_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_17_upstream;
  --niosII_system_burst_17_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_17_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_17_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_17_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_17_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_17_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_17_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_17_upstream_allgrants <= niosII_system_burst_17_upstream_grant_vector;
  --niosII_system_burst_17_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_17_upstream_end_xfer <= NOT ((niosII_system_burst_17_upstream_waits_for_read OR niosII_system_burst_17_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_17_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_17_upstream <= niosII_system_burst_17_upstream_end_xfer AND (((NOT niosII_system_burst_17_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_17_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_17_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_17_upstream AND niosII_system_burst_17_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_17_upstream AND NOT niosII_system_burst_17_upstream_non_bursting_master_requests));
  --niosII_system_burst_17_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_17_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_17_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_17_upstream_arb_share_counter <= niosII_system_burst_17_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_17_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_17_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_17_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_17_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_17_upstream AND NOT niosII_system_burst_17_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_17_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_17_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_17/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_17_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_17_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_17_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_17_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_17/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_17_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_17_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_17_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_17_upstream <= internal_cpu_data_master_requests_niosII_system_burst_17_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_17_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_17_upstream_move_on_to_next_transaction <= niosII_system_burst_17_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_17_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_17_upstream, which is an e_mux
  niosII_system_burst_17_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_17_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_17_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_17_upstream : burstcount_fifo_for_niosII_system_burst_17_upstream_module
    port map(
      data_out => niosII_system_burst_17_upstream_transaction_burst_count,
      empty => niosII_system_burst_17_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input54,
      clk => clk,
      data_in => niosII_system_burst_17_upstream_selected_burstcount,
      read => niosII_system_burst_17_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input55,
      write => module_input56
    );

  module_input54 <= std_logic'('0');
  module_input55 <= std_logic'('0');
  module_input56 <= ((in_a_read_cycle AND NOT niosII_system_burst_17_upstream_waits_for_read) AND niosII_system_burst_17_upstream_load_fifo) AND NOT ((niosII_system_burst_17_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_17_upstream_burstcount_fifo_empty));

  --niosII_system_burst_17_upstream current burst minus one, which is an e_assign
  niosII_system_burst_17_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_17_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_17_upstream, which is an e_mux
  niosII_system_burst_17_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_17_upstream_waits_for_read)) AND NOT niosII_system_burst_17_upstream_load_fifo))) = '1'), niosII_system_burst_17_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_17_upstream_waits_for_read) AND niosII_system_burst_17_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_17_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_17_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_17_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_17_upstream_transaction_burst_count, niosII_system_burst_17_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_17_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_17_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_17_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_17_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_17_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_17_upstream_current_burst <= niosII_system_burst_17_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_17_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_17_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_17_upstream_waits_for_read)) AND niosII_system_burst_17_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_17_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_17_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_17_upstream_waits_for_read)) AND NOT niosII_system_burst_17_upstream_load_fifo) OR niosII_system_burst_17_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_17_upstream_load_fifo <= p0_niosII_system_burst_17_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_17_upstream, which is an e_assign
  niosII_system_burst_17_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_17_upstream_current_burst_minus_one)) AND niosII_system_burst_17_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_17_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_17_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_17_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_17_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_17_upstream,
      full => open,
      clear_fifo => module_input57,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_17_upstream,
      read => niosII_system_burst_17_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input58,
      write => module_input59
    );

  module_input57 <= std_logic'('0');
  module_input58 <= std_logic'('0');
  module_input59 <= in_a_read_cycle AND NOT niosII_system_burst_17_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_17_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_17_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_17_upstream <= niosII_system_burst_17_upstream_readdatavalid_from_sa;
  --niosII_system_burst_17_upstream_writedata mux, which is an e_mux
  niosII_system_burst_17_upstream_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --byteaddress mux for niosII_system_burst_17/upstream, which is an e_mux
  niosII_system_burst_17_upstream_byteaddress <= cpu_data_master_address_to_slave (4 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_17_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_17_upstream;
  --cpu/data_master saved-grant niosII_system_burst_17/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_17_upstream <= internal_cpu_data_master_requests_niosII_system_burst_17_upstream;
  --allow new arb cycle for niosII_system_burst_17/upstream, which is an e_assign
  niosII_system_burst_17_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_17_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_17_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_17_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_17_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_17_upstream_begins_xfer) = '1'), niosII_system_burst_17_upstream_unreg_firsttransfer, niosII_system_burst_17_upstream_reg_firsttransfer);
  --niosII_system_burst_17_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_17_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_17_upstream_slavearbiterlockenable AND niosII_system_burst_17_upstream_any_continuerequest));
  --niosII_system_burst_17_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_17_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_17_upstream_begins_xfer) = '1' then 
        niosII_system_burst_17_upstream_reg_firsttransfer <= niosII_system_burst_17_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_17_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_17_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_17_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_17_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_17_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_17_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_17_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_17_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_17_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_17_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_17_upstream_begins_xfer) = '1' then 
        niosII_system_burst_17_upstream_bbt_burstcounter <= niosII_system_burst_17_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_17_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_17_upstream_beginbursttransfer_internal <= niosII_system_burst_17_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_17_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_17_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_17_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_17_upstream AND cpu_data_master_read;
  --niosII_system_burst_17_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_17_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_17_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_17_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_17_upstream_address mux, which is an e_mux
  niosII_system_burst_17_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_17_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --d1_niosII_system_burst_17_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_17_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_17_upstream_end_xfer <= niosII_system_burst_17_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_17_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_17_upstream_waits_for_read <= niosII_system_burst_17_upstream_in_a_read_cycle AND internal_niosII_system_burst_17_upstream_waitrequest_from_sa;
  --niosII_system_burst_17_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_17_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_17_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_17_upstream_in_a_read_cycle;
  --niosII_system_burst_17_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_17_upstream_waits_for_write <= niosII_system_burst_17_upstream_in_a_write_cycle AND internal_niosII_system_burst_17_upstream_waitrequest_from_sa;
  --niosII_system_burst_17_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_17_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_17_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_17_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_17_upstream_counter <= std_logic'('0');
  --niosII_system_burst_17_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_17_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_17_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_17_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_17_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_17_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_17_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_17_upstream <= internal_cpu_data_master_granted_niosII_system_burst_17_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_17_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_17_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_17_upstream <= internal_cpu_data_master_requests_niosII_system_burst_17_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_17_upstream_burstcount <= internal_niosII_system_burst_17_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_17_upstream_read <= internal_niosII_system_burst_17_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_17_upstream_waitrequest_from_sa <= internal_niosII_system_burst_17_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_17_upstream_write <= internal_niosII_system_burst_17_upstream_write;
--synthesis translate_off
    --niosII_system_burst_17/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line94 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_17_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line94, now);
          write(write_line94, string'(": "));
          write(write_line94, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_17/upstream"));
          write(output, write_line94.all);
          deallocate (write_line94);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_17_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_uart_0_s1_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_17_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_17_downstream_granted_uart_0_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_qualified_request_uart_0_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_read_data_valid_uart_0_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_requests_uart_0_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal uart_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal niosII_system_burst_17_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_17_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_17_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_17_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_17_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_17_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_17_downstream_arbitrator;


architecture europa of niosII_system_burst_17_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_17_downstream_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_17_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_17_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_flush_niosII_system_burst_17_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_17_downstream_qualified_request_uart_0_s1 OR NOT niosII_system_burst_17_downstream_requests_uart_0_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_17_downstream_qualified_request_uart_0_s1 OR NOT ((niosII_system_burst_17_downstream_read OR niosII_system_burst_17_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_uart_0_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_17_downstream_read OR niosII_system_burst_17_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_17_downstream_qualified_request_uart_0_s1 OR NOT ((niosII_system_burst_17_downstream_read OR niosII_system_burst_17_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_uart_0_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_17_downstream_read OR niosII_system_burst_17_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_17_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_17_downstream_address_to_slave <= niosII_system_burst_17_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_17_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_17_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_17_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_17_downstream_read_data_valid_uart_0_s1)))));
  --niosII_system_burst_17/downstream readdata mux, which is an e_mux
  niosII_system_burst_17_downstream_readdata <= uart_0_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_17_downstream_waitrequest <= NOT niosII_system_burst_17_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_17_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_17_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_17_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_17_downstream_address_to_slave <= internal_niosII_system_burst_17_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_17_downstream_waitrequest <= internal_niosII_system_burst_17_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_17_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_17_downstream_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_17_downstream_address_last_time <= niosII_system_burst_17_downstream_address;
      end if;

    end process;

    --niosII_system_burst_17/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_17_downstream_waitrequest AND ((niosII_system_burst_17_downstream_read OR niosII_system_burst_17_downstream_write));
      end if;

    end process;

    --niosII_system_burst_17_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line95 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_17_downstream_address /= niosII_system_burst_17_downstream_address_last_time))))) = '1' then 
          write(write_line95, now);
          write(write_line95, string'(": "));
          write(write_line95, string'("niosII_system_burst_17_downstream_address did not heed wait!!!"));
          write(output, write_line95.all);
          deallocate (write_line95);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_17_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_17_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_17_downstream_burstcount_last_time <= niosII_system_burst_17_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_17_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line96 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_17_downstream_burstcount) /= std_logic'(niosII_system_burst_17_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line96, now);
          write(write_line96, string'(": "));
          write(write_line96, string'("niosII_system_burst_17_downstream_burstcount did not heed wait!!!"));
          write(output, write_line96.all);
          deallocate (write_line96);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_17_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_17_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_17_downstream_byteenable_last_time <= niosII_system_burst_17_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_17_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line97 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_17_downstream_byteenable /= niosII_system_burst_17_downstream_byteenable_last_time))))) = '1' then 
          write(write_line97, now);
          write(write_line97, string'(": "));
          write(write_line97, string'("niosII_system_burst_17_downstream_byteenable did not heed wait!!!"));
          write(output, write_line97.all);
          deallocate (write_line97);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_17_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_17_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_17_downstream_read_last_time <= niosII_system_burst_17_downstream_read;
      end if;

    end process;

    --niosII_system_burst_17_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line98 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_17_downstream_read) /= std_logic'(niosII_system_burst_17_downstream_read_last_time)))))) = '1' then 
          write(write_line98, now);
          write(write_line98, string'(": "));
          write(write_line98, string'("niosII_system_burst_17_downstream_read did not heed wait!!!"));
          write(output, write_line98.all);
          deallocate (write_line98);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_17_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_17_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_17_downstream_write_last_time <= niosII_system_burst_17_downstream_write;
      end if;

    end process;

    --niosII_system_burst_17_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line99 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_17_downstream_write) /= std_logic'(niosII_system_burst_17_downstream_write_last_time)))))) = '1' then 
          write(write_line99, now);
          write(write_line99, string'(": "));
          write(write_line99, string'("niosII_system_burst_17_downstream_write did not heed wait!!!"));
          write(output, write_line99.all);
          deallocate (write_line99);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_17_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_17_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_17_downstream_writedata_last_time <= niosII_system_burst_17_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_17_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line100 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_17_downstream_writedata /= niosII_system_burst_17_downstream_writedata_last_time)))) AND niosII_system_burst_17_downstream_write)) = '1' then 
          write(write_line100, now);
          write(write_line100, string'(": "));
          write(write_line100, string'("niosII_system_burst_17_downstream_writedata did not heed wait!!!"));
          write(output, write_line100.all);
          deallocate (write_line100);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_18_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_18_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_18_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_18_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_18_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_18_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_18_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_18_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_18_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_18_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_18_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_18_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_18_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_18_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_18_upstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_18_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_18_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_18_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_18_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_18_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_18_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_18_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_18_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_18_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity niosII_system_burst_18_upstream_arbitrator;


architecture europa of niosII_system_burst_18_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_18_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_18_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_18_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_18_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_18_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_18_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_18_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_18_upstream_write :  STD_LOGIC;
                signal module_input60 :  STD_LOGIC;
                signal module_input61 :  STD_LOGIC;
                signal module_input62 :  STD_LOGIC;
                signal module_input63 :  STD_LOGIC;
                signal module_input64 :  STD_LOGIC;
                signal module_input65 :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_18_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_18_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_18_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_18_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_18_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_18_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_18_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_18_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_18_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_18_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_18_upstream);
  --assign niosII_system_burst_18_upstream_readdatavalid_from_sa = niosII_system_burst_18_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_18_upstream_readdatavalid_from_sa <= niosII_system_burst_18_upstream_readdatavalid;
  --assign niosII_system_burst_18_upstream_readdata_from_sa = niosII_system_burst_18_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_18_upstream_readdata_from_sa <= niosII_system_burst_18_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_18_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1100100001001000001100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_18_upstream_waitrequest_from_sa = niosII_system_burst_18_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_18_upstream_waitrequest_from_sa <= niosII_system_burst_18_upstream_waitrequest;
  --niosII_system_burst_18_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_18_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_18_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_18_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_18_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_18_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_18_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_18_upstream;
  --niosII_system_burst_18_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_18_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_18_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_18_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_18_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_18_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_18_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_18_upstream_allgrants <= niosII_system_burst_18_upstream_grant_vector;
  --niosII_system_burst_18_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_18_upstream_end_xfer <= NOT ((niosII_system_burst_18_upstream_waits_for_read OR niosII_system_burst_18_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_18_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_18_upstream <= niosII_system_burst_18_upstream_end_xfer AND (((NOT niosII_system_burst_18_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_18_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_18_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_18_upstream AND niosII_system_burst_18_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_18_upstream AND NOT niosII_system_burst_18_upstream_non_bursting_master_requests));
  --niosII_system_burst_18_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_18_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_18_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_18_upstream_arb_share_counter <= niosII_system_burst_18_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_18_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_18_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_18_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_18_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_18_upstream AND NOT niosII_system_burst_18_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_18_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_18_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_18/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_18_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_18_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_18_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_18_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_18/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_18_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_18_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_18_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_18_upstream <= internal_cpu_data_master_requests_niosII_system_burst_18_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_18_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_18_upstream_move_on_to_next_transaction <= niosII_system_burst_18_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_18_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_18_upstream, which is an e_mux
  niosII_system_burst_18_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_18_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_18_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_18_upstream : burstcount_fifo_for_niosII_system_burst_18_upstream_module
    port map(
      data_out => niosII_system_burst_18_upstream_transaction_burst_count,
      empty => niosII_system_burst_18_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input60,
      clk => clk,
      data_in => niosII_system_burst_18_upstream_selected_burstcount,
      read => niosII_system_burst_18_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input61,
      write => module_input62
    );

  module_input60 <= std_logic'('0');
  module_input61 <= std_logic'('0');
  module_input62 <= ((in_a_read_cycle AND NOT niosII_system_burst_18_upstream_waits_for_read) AND niosII_system_burst_18_upstream_load_fifo) AND NOT ((niosII_system_burst_18_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_18_upstream_burstcount_fifo_empty));

  --niosII_system_burst_18_upstream current burst minus one, which is an e_assign
  niosII_system_burst_18_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_18_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_18_upstream, which is an e_mux
  niosII_system_burst_18_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_18_upstream_waits_for_read)) AND NOT niosII_system_burst_18_upstream_load_fifo))) = '1'), niosII_system_burst_18_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_18_upstream_waits_for_read) AND niosII_system_burst_18_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_18_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_18_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_18_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_18_upstream_transaction_burst_count, niosII_system_burst_18_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_18_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_18_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_18_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_18_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_18_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_18_upstream_current_burst <= niosII_system_burst_18_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_18_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_18_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_18_upstream_waits_for_read)) AND niosII_system_burst_18_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_18_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_18_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_18_upstream_waits_for_read)) AND NOT niosII_system_burst_18_upstream_load_fifo) OR niosII_system_burst_18_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_18_upstream_load_fifo <= p0_niosII_system_burst_18_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_18_upstream, which is an e_assign
  niosII_system_burst_18_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_18_upstream_current_burst_minus_one)) AND niosII_system_burst_18_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_18_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_18_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_18_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_18_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_18_upstream,
      full => open,
      clear_fifo => module_input63,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_18_upstream,
      read => niosII_system_burst_18_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input64,
      write => module_input65
    );

  module_input63 <= std_logic'('0');
  module_input64 <= std_logic'('0');
  module_input65 <= in_a_read_cycle AND NOT niosII_system_burst_18_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_18_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_18_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_18_upstream <= niosII_system_burst_18_upstream_readdatavalid_from_sa;
  --niosII_system_burst_18_upstream_writedata mux, which is an e_mux
  niosII_system_burst_18_upstream_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --byteaddress mux for niosII_system_burst_18/upstream, which is an e_mux
  niosII_system_burst_18_upstream_byteaddress <= cpu_data_master_address_to_slave (4 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_18_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_18_upstream;
  --cpu/data_master saved-grant niosII_system_burst_18/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_18_upstream <= internal_cpu_data_master_requests_niosII_system_burst_18_upstream;
  --allow new arb cycle for niosII_system_burst_18/upstream, which is an e_assign
  niosII_system_burst_18_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_18_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_18_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_18_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_18_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_18_upstream_begins_xfer) = '1'), niosII_system_burst_18_upstream_unreg_firsttransfer, niosII_system_burst_18_upstream_reg_firsttransfer);
  --niosII_system_burst_18_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_18_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_18_upstream_slavearbiterlockenable AND niosII_system_burst_18_upstream_any_continuerequest));
  --niosII_system_burst_18_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_18_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_18_upstream_begins_xfer) = '1' then 
        niosII_system_burst_18_upstream_reg_firsttransfer <= niosII_system_burst_18_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_18_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_18_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_18_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_18_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_18_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_18_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_18_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_18_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_18_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_18_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_18_upstream_begins_xfer) = '1' then 
        niosII_system_burst_18_upstream_bbt_burstcounter <= niosII_system_burst_18_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_18_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_18_upstream_beginbursttransfer_internal <= niosII_system_burst_18_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_18_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_18_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_18_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_18_upstream AND cpu_data_master_read;
  --niosII_system_burst_18_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_18_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_18_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_18_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_18_upstream_address mux, which is an e_mux
  niosII_system_burst_18_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_18_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --d1_niosII_system_burst_18_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_18_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_18_upstream_end_xfer <= niosII_system_burst_18_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_18_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_18_upstream_waits_for_read <= niosII_system_burst_18_upstream_in_a_read_cycle AND internal_niosII_system_burst_18_upstream_waitrequest_from_sa;
  --niosII_system_burst_18_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_18_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_18_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_18_upstream_in_a_read_cycle;
  --niosII_system_burst_18_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_18_upstream_waits_for_write <= niosII_system_burst_18_upstream_in_a_write_cycle AND internal_niosII_system_burst_18_upstream_waitrequest_from_sa;
  --niosII_system_burst_18_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_18_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_18_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_18_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_18_upstream_counter <= std_logic'('0');
  --niosII_system_burst_18_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_18_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_18_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_18_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_18_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_18_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_18_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_18_upstream <= internal_cpu_data_master_granted_niosII_system_burst_18_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_18_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_18_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_18_upstream <= internal_cpu_data_master_requests_niosII_system_burst_18_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_18_upstream_burstcount <= internal_niosII_system_burst_18_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_18_upstream_read <= internal_niosII_system_burst_18_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_18_upstream_waitrequest_from_sa <= internal_niosII_system_burst_18_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_18_upstream_write <= internal_niosII_system_burst_18_upstream_write;
--synthesis translate_off
    --niosII_system_burst_18/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line101 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_18_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line101, now);
          write(write_line101, string'(": "));
          write(write_line101, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_18/upstream"));
          write(output, write_line101.all);
          deallocate (write_line101);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_18_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_uart_1_s1_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_18_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_18_downstream_granted_uart_1_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_qualified_request_uart_1_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_read_data_valid_uart_1_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_requests_uart_1_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal uart_1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal niosII_system_burst_18_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_18_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_18_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_18_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_18_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_18_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_18_downstream_arbitrator;


architecture europa of niosII_system_burst_18_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_18_downstream_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_18_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_18_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_flush_niosII_system_burst_18_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_18_downstream_qualified_request_uart_1_s1 OR NOT niosII_system_burst_18_downstream_requests_uart_1_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_18_downstream_qualified_request_uart_1_s1 OR NOT ((niosII_system_burst_18_downstream_read OR niosII_system_burst_18_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_uart_1_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_18_downstream_read OR niosII_system_burst_18_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_18_downstream_qualified_request_uart_1_s1 OR NOT ((niosII_system_burst_18_downstream_read OR niosII_system_burst_18_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_uart_1_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_18_downstream_read OR niosII_system_burst_18_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_18_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_18_downstream_address_to_slave <= niosII_system_burst_18_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_18_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_18_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_18_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_18_downstream_read_data_valid_uart_1_s1)))));
  --niosII_system_burst_18/downstream readdata mux, which is an e_mux
  niosII_system_burst_18_downstream_readdata <= uart_1_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_18_downstream_waitrequest <= NOT niosII_system_burst_18_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_18_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_18_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_18_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_18_downstream_address_to_slave <= internal_niosII_system_burst_18_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_18_downstream_waitrequest <= internal_niosII_system_burst_18_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_18_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_18_downstream_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_18_downstream_address_last_time <= niosII_system_burst_18_downstream_address;
      end if;

    end process;

    --niosII_system_burst_18/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_18_downstream_waitrequest AND ((niosII_system_burst_18_downstream_read OR niosII_system_burst_18_downstream_write));
      end if;

    end process;

    --niosII_system_burst_18_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line102 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_18_downstream_address /= niosII_system_burst_18_downstream_address_last_time))))) = '1' then 
          write(write_line102, now);
          write(write_line102, string'(": "));
          write(write_line102, string'("niosII_system_burst_18_downstream_address did not heed wait!!!"));
          write(output, write_line102.all);
          deallocate (write_line102);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_18_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_18_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_18_downstream_burstcount_last_time <= niosII_system_burst_18_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_18_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line103 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_18_downstream_burstcount) /= std_logic'(niosII_system_burst_18_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line103, now);
          write(write_line103, string'(": "));
          write(write_line103, string'("niosII_system_burst_18_downstream_burstcount did not heed wait!!!"));
          write(output, write_line103.all);
          deallocate (write_line103);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_18_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_18_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_18_downstream_byteenable_last_time <= niosII_system_burst_18_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_18_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line104 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_18_downstream_byteenable /= niosII_system_burst_18_downstream_byteenable_last_time))))) = '1' then 
          write(write_line104, now);
          write(write_line104, string'(": "));
          write(write_line104, string'("niosII_system_burst_18_downstream_byteenable did not heed wait!!!"));
          write(output, write_line104.all);
          deallocate (write_line104);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_18_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_18_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_18_downstream_read_last_time <= niosII_system_burst_18_downstream_read;
      end if;

    end process;

    --niosII_system_burst_18_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line105 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_18_downstream_read) /= std_logic'(niosII_system_burst_18_downstream_read_last_time)))))) = '1' then 
          write(write_line105, now);
          write(write_line105, string'(": "));
          write(write_line105, string'("niosII_system_burst_18_downstream_read did not heed wait!!!"));
          write(output, write_line105.all);
          deallocate (write_line105);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_18_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_18_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_18_downstream_write_last_time <= niosII_system_burst_18_downstream_write;
      end if;

    end process;

    --niosII_system_burst_18_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line106 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_18_downstream_write) /= std_logic'(niosII_system_burst_18_downstream_write_last_time)))))) = '1' then 
          write(write_line106, now);
          write(write_line106, string'(": "));
          write(write_line106, string'("niosII_system_burst_18_downstream_write did not heed wait!!!"));
          write(output, write_line106.all);
          deallocate (write_line106);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_18_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_18_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_18_downstream_writedata_last_time <= niosII_system_burst_18_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_18_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line107 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_18_downstream_writedata /= niosII_system_burst_18_downstream_writedata_last_time)))) AND niosII_system_burst_18_downstream_write)) = '1' then 
          write(write_line107, now);
          write(write_line107, string'(": "));
          write(write_line107, string'("niosII_system_burst_18_downstream_writedata did not heed wait!!!"));
          write(output, write_line107.all);
          deallocate (write_line107);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_19_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_19_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_19_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("00000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("00000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("00000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("00000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_19_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_19_upstream_module;


architecture europa of rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_19_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_19_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : IN STD_LOGIC;
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : IN STD_LOGIC;
                 signal niosII_system_burst_19_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_19_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_19_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_instruction_master_granted_niosII_system_burst_19_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_instruction_master_requests_niosII_system_burst_19_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_19_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_19_upstream_address : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal niosII_system_burst_19_upstream_byteaddress : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
                 signal niosII_system_burst_19_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_19_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_19_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_19_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_19_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_19_upstream_write : OUT STD_LOGIC
              );
end entity niosII_system_burst_19_upstream_arbitrator;


architecture europa of niosII_system_burst_19_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_19_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_19_upstream_module;

component rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_19_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_19_upstream_module;

                signal cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_output_from_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal cpu_instruction_master_saved_grant_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_instruction_master_granted_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal internal_cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal internal_cpu_instruction_master_requests_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_19_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal module_input66 :  STD_LOGIC;
                signal module_input67 :  STD_LOGIC;
                signal module_input68 :  STD_LOGIC;
                signal module_input69 :  STD_LOGIC;
                signal module_input70 :  STD_LOGIC;
                signal module_input71 :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_19_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_19_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_19_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_current_burst :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_19_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_19_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_next_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_19_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_selected_burstcount :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_19_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_19_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_19_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_19_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_19_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_19_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream);
  --assign niosII_system_burst_19_upstream_readdatavalid_from_sa = niosII_system_burst_19_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_19_upstream_readdatavalid_from_sa <= niosII_system_burst_19_upstream_readdatavalid;
  --assign niosII_system_burst_19_upstream_readdata_from_sa = niosII_system_burst_19_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_19_upstream_readdata_from_sa <= niosII_system_burst_19_upstream_readdata;
  internal_cpu_instruction_master_requests_niosII_system_burst_19_upstream <= ((to_std_logic(((Std_Logic_Vector'(cpu_instruction_master_address_to_slave(24 DOWNTO 19) & std_logic_vector'("0000000000000000000")) = std_logic_vector'("1100010000000000000000000")))) AND (cpu_instruction_master_read))) AND cpu_instruction_master_read;
  --assign niosII_system_burst_19_upstream_waitrequest_from_sa = niosII_system_burst_19_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_19_upstream_waitrequest_from_sa <= niosII_system_burst_19_upstream_waitrequest;
  --niosII_system_burst_19_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_19_upstream_arb_share_set_values <= std_logic_vector'("00000001");
  --niosII_system_burst_19_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_19_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_19_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_19_upstream_any_bursting_master_saved_grant <= cpu_instruction_master_saved_grant_niosII_system_burst_19_upstream;
  --niosII_system_burst_19_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_19_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_19_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_19_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_19_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_19_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_19_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_19_upstream_allgrants <= niosII_system_burst_19_upstream_grant_vector;
  --niosII_system_burst_19_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_19_upstream_end_xfer <= NOT ((niosII_system_burst_19_upstream_waits_for_read OR niosII_system_burst_19_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_19_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_19_upstream <= niosII_system_burst_19_upstream_end_xfer AND (((NOT niosII_system_burst_19_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_19_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_19_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_19_upstream AND niosII_system_burst_19_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_19_upstream AND NOT niosII_system_burst_19_upstream_non_bursting_master_requests));
  --niosII_system_burst_19_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_19_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_19_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_19_upstream_arb_share_counter <= niosII_system_burst_19_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_19_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_19_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_19_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_19_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_19_upstream AND NOT niosII_system_burst_19_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_19_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_19_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/instruction_master niosII_system_burst_19/upstream arbiterlock, which is an e_assign
  cpu_instruction_master_arbiterlock <= niosII_system_burst_19_upstream_slavearbiterlockenable AND cpu_instruction_master_continuerequest;
  --niosII_system_burst_19_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_19_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_19_upstream_arb_share_counter_next_value);
  --cpu/instruction_master niosII_system_burst_19/upstream arbiterlock2, which is an e_assign
  cpu_instruction_master_arbiterlock2 <= niosII_system_burst_19_upstream_slavearbiterlockenable2 AND cpu_instruction_master_continuerequest;
  --niosII_system_burst_19_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_19_upstream_any_continuerequest <= std_logic'('1');
  --cpu_instruction_master_continuerequest continued request, which is an e_assign
  cpu_instruction_master_continuerequest <= std_logic'('1');
  internal_cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_19_upstream AND NOT ((cpu_instruction_master_read AND (((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_latency_counter))))))) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register)))));
  --unique name for niosII_system_burst_19_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_19_upstream_move_on_to_next_transaction <= niosII_system_burst_19_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_19_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_19_upstream, which is an e_mux
  niosII_system_burst_19_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_niosII_system_burst_19_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_instruction_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --burstcount_fifo_for_niosII_system_burst_19_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_19_upstream : burstcount_fifo_for_niosII_system_burst_19_upstream_module
    port map(
      data_out => niosII_system_burst_19_upstream_transaction_burst_count,
      empty => niosII_system_burst_19_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input66,
      clk => clk,
      data_in => niosII_system_burst_19_upstream_selected_burstcount,
      read => niosII_system_burst_19_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input67,
      write => module_input68
    );

  module_input66 <= std_logic'('0');
  module_input67 <= std_logic'('0');
  module_input68 <= ((in_a_read_cycle AND NOT niosII_system_burst_19_upstream_waits_for_read) AND niosII_system_burst_19_upstream_load_fifo) AND NOT ((niosII_system_burst_19_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_19_upstream_burstcount_fifo_empty));

  --niosII_system_burst_19_upstream current burst minus one, which is an e_assign
  niosII_system_burst_19_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_19_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --what to load in current_burst, for niosII_system_burst_19_upstream, which is an e_mux
  niosII_system_burst_19_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_19_upstream_waits_for_read)) AND NOT niosII_system_burst_19_upstream_load_fifo))) = '1'), (niosII_system_burst_19_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_19_upstream_waits_for_read) AND niosII_system_burst_19_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_19_upstream_burstcount_fifo_empty))) = '1'), (niosII_system_burst_19_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'((niosII_system_burst_19_upstream_this_cycle_is_the_last_burst)) = '1'), (niosII_system_burst_19_upstream_transaction_burst_count & A_ToStdLogicVector(std_logic'('0'))), (std_logic_vector'("0") & (niosII_system_burst_19_upstream_current_burst_minus_one))))), 5);
  --the current burst count for niosII_system_burst_19_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_19_upstream_current_burst <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_19_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_19_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_19_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_19_upstream_current_burst <= niosII_system_burst_19_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_19_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_19_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_19_upstream_waits_for_read)) AND niosII_system_burst_19_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_19_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_19_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_19_upstream_waits_for_read)) AND NOT niosII_system_burst_19_upstream_load_fifo) OR niosII_system_burst_19_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_19_upstream_load_fifo <= p0_niosII_system_burst_19_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_19_upstream, which is an e_assign
  niosII_system_burst_19_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_19_upstream_current_burst_minus_one)) AND niosII_system_burst_19_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_19_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_19_upstream : rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_19_upstream_module
    port map(
      data_out => cpu_instruction_master_rdv_fifo_output_from_niosII_system_burst_19_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_19_upstream,
      full => open,
      clear_fifo => module_input69,
      clk => clk,
      data_in => internal_cpu_instruction_master_granted_niosII_system_burst_19_upstream,
      read => niosII_system_burst_19_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input70,
      write => module_input71
    );

  module_input69 <= std_logic'('0');
  module_input70 <= std_logic'('0');
  module_input71 <= in_a_read_cycle AND NOT niosII_system_burst_19_upstream_waits_for_read;

  cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register <= NOT cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_19_upstream;
  --local readdatavalid cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream, which is an e_mux
  cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream <= niosII_system_burst_19_upstream_readdatavalid_from_sa;
  --byteaddress mux for niosII_system_burst_19/upstream, which is an e_mux
  niosII_system_burst_19_upstream_byteaddress <= cpu_instruction_master_address_to_slave (19 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_instruction_master_granted_niosII_system_burst_19_upstream <= internal_cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream;
  --cpu/instruction_master saved-grant niosII_system_burst_19/upstream, which is an e_assign
  cpu_instruction_master_saved_grant_niosII_system_burst_19_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_19_upstream;
  --allow new arb cycle for niosII_system_burst_19/upstream, which is an e_assign
  niosII_system_burst_19_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_19_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_19_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_19_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_19_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_19_upstream_begins_xfer) = '1'), niosII_system_burst_19_upstream_unreg_firsttransfer, niosII_system_burst_19_upstream_reg_firsttransfer);
  --niosII_system_burst_19_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_19_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_19_upstream_slavearbiterlockenable AND niosII_system_burst_19_upstream_any_continuerequest));
  --niosII_system_burst_19_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_19_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_19_upstream_begins_xfer) = '1' then 
        niosII_system_burst_19_upstream_reg_firsttransfer <= niosII_system_burst_19_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_19_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_19_upstream_beginbursttransfer_internal <= niosII_system_burst_19_upstream_begins_xfer;
  --niosII_system_burst_19_upstream_read assignment, which is an e_mux
  niosII_system_burst_19_upstream_read <= internal_cpu_instruction_master_granted_niosII_system_burst_19_upstream AND cpu_instruction_master_read;
  --niosII_system_burst_19_upstream_write assignment, which is an e_mux
  niosII_system_burst_19_upstream_write <= std_logic'('0');
  --niosII_system_burst_19_upstream_address mux, which is an e_mux
  niosII_system_burst_19_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(cpu_instruction_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 19);
  --d1_niosII_system_burst_19_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_19_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_19_upstream_end_xfer <= niosII_system_burst_19_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_19_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_19_upstream_waits_for_read <= niosII_system_burst_19_upstream_in_a_read_cycle AND internal_niosII_system_burst_19_upstream_waitrequest_from_sa;
  --niosII_system_burst_19_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_19_upstream_in_a_read_cycle <= internal_cpu_instruction_master_granted_niosII_system_burst_19_upstream AND cpu_instruction_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_19_upstream_in_a_read_cycle;
  --niosII_system_burst_19_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_19_upstream_waits_for_write <= niosII_system_burst_19_upstream_in_a_write_cycle AND internal_niosII_system_burst_19_upstream_waitrequest_from_sa;
  --niosII_system_burst_19_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_19_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_19_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_19_upstream_counter <= std_logic'('0');
  --niosII_system_burst_19_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_19_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 2);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_19_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_instruction_master_granted_niosII_system_burst_19_upstream <= internal_cpu_instruction_master_granted_niosII_system_burst_19_upstream;
  --vhdl renameroo for output signals
  cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream <= internal_cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream;
  --vhdl renameroo for output signals
  cpu_instruction_master_requests_niosII_system_burst_19_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_19_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_19_upstream_waitrequest_from_sa <= internal_niosII_system_burst_19_upstream_waitrequest_from_sa;
--synthesis translate_off
    --niosII_system_burst_19/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/instruction_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line108 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_instruction_master_requests_niosII_system_burst_19_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_instruction_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line108, now);
          write(write_line108, string'(": "));
          write(write_line108, string'("cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_19/upstream"));
          write(output, write_line108.all);
          deallocate (write_line108);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_19_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_tsb_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal incoming_sram_IF_0_tsb_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_address : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_granted_sram_IF_0_tsb : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_requests_sram_IF_0_tsb : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_19_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_19_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_19_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_19_downstream_arbitrator;


architecture europa of niosII_system_burst_19_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_19_downstream_address_to_slave :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal internal_niosII_system_burst_19_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_niosII_system_burst_19_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_19_downstream_address_last_time :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_19_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_19_downstream_is_granted_some_slave :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_niosII_system_burst_19_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pre_flush_niosII_system_burst_19_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb OR NOT niosII_system_burst_19_downstream_requests_sram_IF_0_tsb)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_19_downstream_granted_sram_IF_0_tsb OR NOT niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb OR NOT niosII_system_burst_19_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_tsb_avalon_slave_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_19_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb OR NOT niosII_system_burst_19_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_19_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_19_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_19_downstream_address_to_slave <= niosII_system_burst_19_downstream_address;
  --niosII_system_burst_19_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_19_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_19_downstream_read_but_no_slave_selected <= (niosII_system_burst_19_downstream_read AND niosII_system_burst_19_downstream_run) AND NOT niosII_system_burst_19_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  niosII_system_burst_19_downstream_is_granted_some_slave <= niosII_system_burst_19_downstream_granted_sram_IF_0_tsb;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_19_downstream_readdatavalid <= niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb;
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_19_downstream_readdatavalid <= niosII_system_burst_19_downstream_read_but_no_slave_selected OR pre_flush_niosII_system_burst_19_downstream_readdatavalid;
  --niosII_system_burst_19/downstream readdata mux, which is an e_mux
  niosII_system_burst_19_downstream_readdata <= incoming_sram_IF_0_tsb_data;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_19_downstream_waitrequest <= NOT niosII_system_burst_19_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_niosII_system_burst_19_downstream_latency_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      internal_niosII_system_burst_19_downstream_latency_counter <= p1_niosII_system_burst_19_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_niosII_system_burst_19_downstream_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((niosII_system_burst_19_downstream_run AND niosII_system_burst_19_downstream_read))) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_niosII_system_burst_19_downstream_latency_counter)) /= std_logic_vector'("00")), ((std_logic_vector'("0000000000000000000000000000000") & (internal_niosII_system_burst_19_downstream_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (A_REP(niosII_system_burst_19_downstream_requests_sram_IF_0_tsb, 2))) AND std_logic_vector'("00000000000000000000000000000010")), 2);
  --niosII_system_burst_19_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_19_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_19_downstream_address_to_slave <= internal_niosII_system_burst_19_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_19_downstream_latency_counter <= internal_niosII_system_burst_19_downstream_latency_counter;
  --vhdl renameroo for output signals
  niosII_system_burst_19_downstream_waitrequest <= internal_niosII_system_burst_19_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_19_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_19_downstream_address_last_time <= std_logic_vector'("0000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_19_downstream_address_last_time <= niosII_system_burst_19_downstream_address;
      end if;

    end process;

    --niosII_system_burst_19/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_19_downstream_waitrequest AND ((niosII_system_burst_19_downstream_read OR niosII_system_burst_19_downstream_write));
      end if;

    end process;

    --niosII_system_burst_19_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line109 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_19_downstream_address /= niosII_system_burst_19_downstream_address_last_time))))) = '1' then 
          write(write_line109, now);
          write(write_line109, string'(": "));
          write(write_line109, string'("niosII_system_burst_19_downstream_address did not heed wait!!!"));
          write(output, write_line109.all);
          deallocate (write_line109);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_19_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_19_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_19_downstream_burstcount_last_time <= niosII_system_burst_19_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_19_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line110 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_19_downstream_burstcount) /= std_logic'(niosII_system_burst_19_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line110, now);
          write(write_line110, string'(": "));
          write(write_line110, string'("niosII_system_burst_19_downstream_burstcount did not heed wait!!!"));
          write(output, write_line110.all);
          deallocate (write_line110);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_19_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_19_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_19_downstream_byteenable_last_time <= niosII_system_burst_19_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_19_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line111 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_19_downstream_byteenable /= niosII_system_burst_19_downstream_byteenable_last_time))))) = '1' then 
          write(write_line111, now);
          write(write_line111, string'(": "));
          write(write_line111, string'("niosII_system_burst_19_downstream_byteenable did not heed wait!!!"));
          write(output, write_line111.all);
          deallocate (write_line111);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_19_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_19_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_19_downstream_read_last_time <= niosII_system_burst_19_downstream_read;
      end if;

    end process;

    --niosII_system_burst_19_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line112 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_19_downstream_read) /= std_logic'(niosII_system_burst_19_downstream_read_last_time)))))) = '1' then 
          write(write_line112, now);
          write(write_line112, string'(": "));
          write(write_line112, string'("niosII_system_burst_19_downstream_read did not heed wait!!!"));
          write(output, write_line112.all);
          deallocate (write_line112);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_19_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_19_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_19_downstream_write_last_time <= niosII_system_burst_19_downstream_write;
      end if;

    end process;

    --niosII_system_burst_19_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line113 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_19_downstream_write) /= std_logic'(niosII_system_burst_19_downstream_write_last_time)))))) = '1' then 
          write(write_line113, now);
          write(write_line113, string'(": "));
          write(write_line113, string'("niosII_system_burst_19_downstream_write did not heed wait!!!"));
          write(output, write_line113.all);
          deallocate (write_line113);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_19_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_19_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_19_downstream_writedata_last_time <= niosII_system_burst_19_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_19_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line114 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_19_downstream_writedata /= niosII_system_burst_19_downstream_writedata_last_time)))) AND niosII_system_burst_19_downstream_write)) = '1' then 
          write(write_line114, now);
          write(write_line114, string'(": "));
          write(write_line114, string'("niosII_system_burst_19_downstream_writedata did not heed wait!!!"));
          write(output, write_line114.all);
          deallocate (write_line114);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_2_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_2_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_2_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("0000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_2_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_2_upstream_module;


architecture europa of rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_2_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_2_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : IN STD_LOGIC;
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : IN STD_LOGIC;
                 signal niosII_system_burst_2_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_2_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_2_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_instruction_master_granted_niosII_system_burst_2_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_instruction_master_requests_niosII_system_burst_2_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_2_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_2_upstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal niosII_system_burst_2_upstream_byteaddress : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_2_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_2_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_2_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_2_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_2_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_2_upstream_write : OUT STD_LOGIC
              );
end entity niosII_system_burst_2_upstream_arbitrator;


architecture europa of niosII_system_burst_2_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_2_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_2_upstream_module;

component rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_2_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_2_upstream_module;

                signal cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_output_from_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal cpu_instruction_master_saved_grant_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_instruction_master_granted_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal internal_cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal internal_cpu_instruction_master_requests_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_2_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal module_input72 :  STD_LOGIC;
                signal module_input73 :  STD_LOGIC;
                signal module_input74 :  STD_LOGIC;
                signal module_input75 :  STD_LOGIC;
                signal module_input76 :  STD_LOGIC;
                signal module_input77 :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_2_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_2_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_2_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_2_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_2_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_2_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_2_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_2_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_2_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_2_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_2_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_2_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream);
  --assign niosII_system_burst_2_upstream_readdatavalid_from_sa = niosII_system_burst_2_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_2_upstream_readdatavalid_from_sa <= niosII_system_burst_2_upstream_readdatavalid;
  --assign niosII_system_burst_2_upstream_readdata_from_sa = niosII_system_burst_2_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_2_upstream_readdata_from_sa <= niosII_system_burst_2_upstream_readdata;
  internal_cpu_instruction_master_requests_niosII_system_burst_2_upstream <= ((to_std_logic(((Std_Logic_Vector'(cpu_instruction_master_address_to_slave(24 DOWNTO 14) & std_logic_vector'("00000000000000")) = std_logic_vector'("1100100000100000000000000")))) AND (cpu_instruction_master_read))) AND cpu_instruction_master_read;
  --assign niosII_system_burst_2_upstream_waitrequest_from_sa = niosII_system_burst_2_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_2_upstream_waitrequest_from_sa <= niosII_system_burst_2_upstream_waitrequest;
  --niosII_system_burst_2_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_2_upstream_arb_share_set_values <= std_logic_vector'("00000001");
  --niosII_system_burst_2_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_2_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_2_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_2_upstream_any_bursting_master_saved_grant <= cpu_instruction_master_saved_grant_niosII_system_burst_2_upstream;
  --niosII_system_burst_2_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_2_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_2_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_2_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_2_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_2_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_2_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_2_upstream_allgrants <= niosII_system_burst_2_upstream_grant_vector;
  --niosII_system_burst_2_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_2_upstream_end_xfer <= NOT ((niosII_system_burst_2_upstream_waits_for_read OR niosII_system_burst_2_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_2_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_2_upstream <= niosII_system_burst_2_upstream_end_xfer AND (((NOT niosII_system_burst_2_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_2_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_2_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_2_upstream AND niosII_system_burst_2_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_2_upstream AND NOT niosII_system_burst_2_upstream_non_bursting_master_requests));
  --niosII_system_burst_2_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_2_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_2_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_2_upstream_arb_share_counter <= niosII_system_burst_2_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_2_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_2_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_2_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_2_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_2_upstream AND NOT niosII_system_burst_2_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_2_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_2_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/instruction_master niosII_system_burst_2/upstream arbiterlock, which is an e_assign
  cpu_instruction_master_arbiterlock <= niosII_system_burst_2_upstream_slavearbiterlockenable AND cpu_instruction_master_continuerequest;
  --niosII_system_burst_2_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_2_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_2_upstream_arb_share_counter_next_value);
  --cpu/instruction_master niosII_system_burst_2/upstream arbiterlock2, which is an e_assign
  cpu_instruction_master_arbiterlock2 <= niosII_system_burst_2_upstream_slavearbiterlockenable2 AND cpu_instruction_master_continuerequest;
  --niosII_system_burst_2_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_2_upstream_any_continuerequest <= std_logic'('1');
  --cpu_instruction_master_continuerequest continued request, which is an e_assign
  cpu_instruction_master_continuerequest <= std_logic'('1');
  internal_cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_2_upstream AND NOT ((cpu_instruction_master_read AND (((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_latency_counter))))))) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register)) OR (cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register)))));
  --unique name for niosII_system_burst_2_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_2_upstream_move_on_to_next_transaction <= niosII_system_burst_2_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_2_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_2_upstream, which is an e_mux
  niosII_system_burst_2_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_niosII_system_burst_2_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_instruction_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_2_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_2_upstream : burstcount_fifo_for_niosII_system_burst_2_upstream_module
    port map(
      data_out => niosII_system_burst_2_upstream_transaction_burst_count,
      empty => niosII_system_burst_2_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input72,
      clk => clk,
      data_in => niosII_system_burst_2_upstream_selected_burstcount,
      read => niosII_system_burst_2_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input73,
      write => module_input74
    );

  module_input72 <= std_logic'('0');
  module_input73 <= std_logic'('0');
  module_input74 <= ((in_a_read_cycle AND NOT niosII_system_burst_2_upstream_waits_for_read) AND niosII_system_burst_2_upstream_load_fifo) AND NOT ((niosII_system_burst_2_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_2_upstream_burstcount_fifo_empty));

  --niosII_system_burst_2_upstream current burst minus one, which is an e_assign
  niosII_system_burst_2_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_2_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_2_upstream, which is an e_mux
  niosII_system_burst_2_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_2_upstream_waits_for_read)) AND NOT niosII_system_burst_2_upstream_load_fifo))) = '1'), niosII_system_burst_2_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_2_upstream_waits_for_read) AND niosII_system_burst_2_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_2_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_2_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_2_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_2_upstream_transaction_burst_count, niosII_system_burst_2_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_2_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_2_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_2_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_2_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_2_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_2_upstream_current_burst <= niosII_system_burst_2_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_2_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_2_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_2_upstream_waits_for_read)) AND niosII_system_burst_2_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_2_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_2_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_2_upstream_waits_for_read)) AND NOT niosII_system_burst_2_upstream_load_fifo) OR niosII_system_burst_2_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_2_upstream_load_fifo <= p0_niosII_system_burst_2_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_2_upstream, which is an e_assign
  niosII_system_burst_2_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_2_upstream_current_burst_minus_one)) AND niosII_system_burst_2_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_2_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_2_upstream : rdv_fifo_for_cpu_instruction_master_to_niosII_system_burst_2_upstream_module
    port map(
      data_out => cpu_instruction_master_rdv_fifo_output_from_niosII_system_burst_2_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_2_upstream,
      full => open,
      clear_fifo => module_input75,
      clk => clk,
      data_in => internal_cpu_instruction_master_granted_niosII_system_burst_2_upstream,
      read => niosII_system_burst_2_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input76,
      write => module_input77
    );

  module_input75 <= std_logic'('0');
  module_input76 <= std_logic'('0');
  module_input77 <= in_a_read_cycle AND NOT niosII_system_burst_2_upstream_waits_for_read;

  cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register <= NOT cpu_instruction_master_rdv_fifo_empty_niosII_system_burst_2_upstream;
  --local readdatavalid cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream, which is an e_mux
  cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream <= niosII_system_burst_2_upstream_readdatavalid_from_sa;
  --byteaddress mux for niosII_system_burst_2/upstream, which is an e_mux
  niosII_system_burst_2_upstream_byteaddress <= cpu_instruction_master_address_to_slave (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_instruction_master_granted_niosII_system_burst_2_upstream <= internal_cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream;
  --cpu/instruction_master saved-grant niosII_system_burst_2/upstream, which is an e_assign
  cpu_instruction_master_saved_grant_niosII_system_burst_2_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_2_upstream;
  --allow new arb cycle for niosII_system_burst_2/upstream, which is an e_assign
  niosII_system_burst_2_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_2_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_2_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_2_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_2_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_2_upstream_begins_xfer) = '1'), niosII_system_burst_2_upstream_unreg_firsttransfer, niosII_system_burst_2_upstream_reg_firsttransfer);
  --niosII_system_burst_2_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_2_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_2_upstream_slavearbiterlockenable AND niosII_system_burst_2_upstream_any_continuerequest));
  --niosII_system_burst_2_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_2_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_2_upstream_begins_xfer) = '1' then 
        niosII_system_burst_2_upstream_reg_firsttransfer <= niosII_system_burst_2_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_2_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_2_upstream_beginbursttransfer_internal <= niosII_system_burst_2_upstream_begins_xfer;
  --niosII_system_burst_2_upstream_read assignment, which is an e_mux
  niosII_system_burst_2_upstream_read <= internal_cpu_instruction_master_granted_niosII_system_burst_2_upstream AND cpu_instruction_master_read;
  --niosII_system_burst_2_upstream_write assignment, which is an e_mux
  niosII_system_burst_2_upstream_write <= std_logic'('0');
  --niosII_system_burst_2_upstream_address mux, which is an e_mux
  niosII_system_burst_2_upstream_address <= cpu_instruction_master_address_to_slave (13 DOWNTO 0);
  --d1_niosII_system_burst_2_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_2_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_2_upstream_end_xfer <= niosII_system_burst_2_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_2_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_2_upstream_waits_for_read <= niosII_system_burst_2_upstream_in_a_read_cycle AND internal_niosII_system_burst_2_upstream_waitrequest_from_sa;
  --niosII_system_burst_2_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_2_upstream_in_a_read_cycle <= internal_cpu_instruction_master_granted_niosII_system_burst_2_upstream AND cpu_instruction_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_2_upstream_in_a_read_cycle;
  --niosII_system_burst_2_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_2_upstream_waits_for_write <= niosII_system_burst_2_upstream_in_a_write_cycle AND internal_niosII_system_burst_2_upstream_waitrequest_from_sa;
  --niosII_system_burst_2_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_2_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_2_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_2_upstream_counter <= std_logic'('0');
  --niosII_system_burst_2_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_2_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_2_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_instruction_master_granted_niosII_system_burst_2_upstream <= internal_cpu_instruction_master_granted_niosII_system_burst_2_upstream;
  --vhdl renameroo for output signals
  cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream <= internal_cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream;
  --vhdl renameroo for output signals
  cpu_instruction_master_requests_niosII_system_burst_2_upstream <= internal_cpu_instruction_master_requests_niosII_system_burst_2_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_2_upstream_waitrequest_from_sa <= internal_niosII_system_burst_2_upstream_waitrequest_from_sa;
--synthesis translate_off
    --niosII_system_burst_2/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/instruction_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line115 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_instruction_master_requests_niosII_system_burst_2_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_instruction_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line115, now);
          write(write_line115, string'(": "));
          write(write_line115, string'("cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_2/upstream"));
          write(output, write_line115.all);
          deallocate (write_line115);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_2_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_memory_s1_end_xfer : IN STD_LOGIC;
                 signal memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_2_downstream_address : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal niosII_system_burst_2_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_2_downstream_granted_memory_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_qualified_request_memory_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_read_data_valid_memory_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_requests_memory_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_2_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal niosII_system_burst_2_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_2_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_2_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_2_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_2_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_2_downstream_arbitrator;


architecture europa of niosII_system_burst_2_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_2_downstream_address_to_slave :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal internal_niosII_system_burst_2_downstream_latency_counter :  STD_LOGIC;
                signal internal_niosII_system_burst_2_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_address_last_time :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_2_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_2_downstream_is_granted_some_slave :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_niosII_system_burst_2_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_niosII_system_burst_2_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_2_downstream_qualified_request_memory_s1 OR NOT niosII_system_burst_2_downstream_requests_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_2_downstream_granted_memory_s1 OR NOT niosII_system_burst_2_downstream_qualified_request_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_2_downstream_qualified_request_memory_s1 OR NOT ((niosII_system_burst_2_downstream_read OR niosII_system_burst_2_downstream_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_2_downstream_read OR niosII_system_burst_2_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_2_downstream_qualified_request_memory_s1 OR NOT ((niosII_system_burst_2_downstream_read OR niosII_system_burst_2_downstream_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_2_downstream_read OR niosII_system_burst_2_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_2_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_2_downstream_address_to_slave <= niosII_system_burst_2_downstream_address;
  --niosII_system_burst_2_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_2_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_2_downstream_read_but_no_slave_selected <= (niosII_system_burst_2_downstream_read AND niosII_system_burst_2_downstream_run) AND NOT niosII_system_burst_2_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  niosII_system_burst_2_downstream_is_granted_some_slave <= niosII_system_burst_2_downstream_granted_memory_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_2_downstream_readdatavalid <= niosII_system_burst_2_downstream_read_data_valid_memory_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_2_downstream_readdatavalid <= niosII_system_burst_2_downstream_read_but_no_slave_selected OR pre_flush_niosII_system_burst_2_downstream_readdatavalid;
  --niosII_system_burst_2/downstream readdata mux, which is an e_mux
  niosII_system_burst_2_downstream_readdata <= memory_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_2_downstream_waitrequest <= NOT niosII_system_burst_2_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_niosII_system_burst_2_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_niosII_system_burst_2_downstream_latency_counter <= p1_niosII_system_burst_2_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_niosII_system_burst_2_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((niosII_system_burst_2_downstream_run AND niosII_system_burst_2_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_2_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_2_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_2_downstream_requests_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --niosII_system_burst_2_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_2_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_2_downstream_address_to_slave <= internal_niosII_system_burst_2_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_2_downstream_latency_counter <= internal_niosII_system_burst_2_downstream_latency_counter;
  --vhdl renameroo for output signals
  niosII_system_burst_2_downstream_waitrequest <= internal_niosII_system_burst_2_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_2_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_2_downstream_address_last_time <= std_logic_vector'("00000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_2_downstream_address_last_time <= niosII_system_burst_2_downstream_address;
      end if;

    end process;

    --niosII_system_burst_2/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_2_downstream_waitrequest AND ((niosII_system_burst_2_downstream_read OR niosII_system_burst_2_downstream_write));
      end if;

    end process;

    --niosII_system_burst_2_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line116 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_2_downstream_address /= niosII_system_burst_2_downstream_address_last_time))))) = '1' then 
          write(write_line116, now);
          write(write_line116, string'(": "));
          write(write_line116, string'("niosII_system_burst_2_downstream_address did not heed wait!!!"));
          write(output, write_line116.all);
          deallocate (write_line116);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_2_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_2_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_2_downstream_burstcount_last_time <= niosII_system_burst_2_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_2_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line117 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_2_downstream_burstcount) /= std_logic'(niosII_system_burst_2_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line117, now);
          write(write_line117, string'(": "));
          write(write_line117, string'("niosII_system_burst_2_downstream_burstcount did not heed wait!!!"));
          write(output, write_line117.all);
          deallocate (write_line117);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_2_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_2_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_2_downstream_byteenable_last_time <= niosII_system_burst_2_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_2_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line118 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_2_downstream_byteenable /= niosII_system_burst_2_downstream_byteenable_last_time))))) = '1' then 
          write(write_line118, now);
          write(write_line118, string'(": "));
          write(write_line118, string'("niosII_system_burst_2_downstream_byteenable did not heed wait!!!"));
          write(output, write_line118.all);
          deallocate (write_line118);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_2_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_2_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_2_downstream_read_last_time <= niosII_system_burst_2_downstream_read;
      end if;

    end process;

    --niosII_system_burst_2_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line119 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_2_downstream_read) /= std_logic'(niosII_system_burst_2_downstream_read_last_time)))))) = '1' then 
          write(write_line119, now);
          write(write_line119, string'(": "));
          write(write_line119, string'("niosII_system_burst_2_downstream_read did not heed wait!!!"));
          write(output, write_line119.all);
          deallocate (write_line119);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_2_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_2_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_2_downstream_write_last_time <= niosII_system_burst_2_downstream_write;
      end if;

    end process;

    --niosII_system_burst_2_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line120 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_2_downstream_write) /= std_logic'(niosII_system_burst_2_downstream_write_last_time)))))) = '1' then 
          write(write_line120, now);
          write(write_line120, string'(": "));
          write(write_line120, string'("niosII_system_burst_2_downstream_write did not heed wait!!!"));
          write(output, write_line120.all);
          deallocate (write_line120);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_2_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_2_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_2_downstream_writedata_last_time <= niosII_system_burst_2_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_2_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line121 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_2_downstream_writedata /= niosII_system_burst_2_downstream_writedata_last_time)))) AND niosII_system_burst_2_downstream_write)) = '1' then 
          write(write_line121, now);
          write(write_line121, string'(": "));
          write(write_line121, string'("niosII_system_burst_2_downstream_writedata did not heed wait!!!"));
          write(output, write_line121.all);
          deallocate (write_line121);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_20_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_20_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_20_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("00000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("00000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("00000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("00000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_20_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_20_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_20_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_20_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal niosII_system_burst_20_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_20_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_20_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_byteenable_niosII_system_burst_20_upstream : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_granted_niosII_system_burst_20_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_20_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_20_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_20_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_20_upstream_address : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal niosII_system_burst_20_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_20_upstream_byteaddress : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
                 signal niosII_system_burst_20_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_20_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_20_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_20_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_20_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_20_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_20_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity niosII_system_burst_20_upstream_arbitrator;


architecture europa of niosII_system_burst_20_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_20_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_20_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_20_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_20_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_byteenable_niosII_system_burst_20_upstream_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_byteenable_niosII_system_burst_20_upstream_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_byteenable_niosII_system_burst_20_upstream :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_data_master_granted_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_20_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_20_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_20_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_20_upstream_write :  STD_LOGIC;
                signal module_input78 :  STD_LOGIC;
                signal module_input79 :  STD_LOGIC;
                signal module_input80 :  STD_LOGIC;
                signal module_input81 :  STD_LOGIC;
                signal module_input82 :  STD_LOGIC;
                signal module_input83 :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_20_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_20_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_20_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_20_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_current_burst :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_20_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_20_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_20_upstream_next_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_20_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_selected_burstcount :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_20_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_20_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_20_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_20_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_20_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_20_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_20_upstream);
  --assign niosII_system_burst_20_upstream_readdatavalid_from_sa = niosII_system_burst_20_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_20_upstream_readdatavalid_from_sa <= niosII_system_burst_20_upstream_readdatavalid;
  --assign niosII_system_burst_20_upstream_readdata_from_sa = niosII_system_burst_20_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_20_upstream_readdata_from_sa <= niosII_system_burst_20_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_20_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 19) & std_logic_vector'("0000000000000000000")) = std_logic_vector'("1100010000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_20_upstream_waitrequest_from_sa = niosII_system_burst_20_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_20_upstream_waitrequest_from_sa <= niosII_system_burst_20_upstream_waitrequest;
  --niosII_system_burst_20_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_20_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_20_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (A_SLL(cpu_data_master_burstcount,std_logic_vector'("00000000000000000000000000000001")))), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_20_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_20_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_20_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_20_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_20_upstream;
  --niosII_system_burst_20_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_20_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_20_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_20_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_20_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_20_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_20_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_20_upstream_allgrants <= niosII_system_burst_20_upstream_grant_vector;
  --niosII_system_burst_20_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_20_upstream_end_xfer <= NOT ((niosII_system_burst_20_upstream_waits_for_read OR niosII_system_burst_20_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_20_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_20_upstream <= niosII_system_burst_20_upstream_end_xfer AND (((NOT niosII_system_burst_20_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_20_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_20_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_20_upstream AND niosII_system_burst_20_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_20_upstream AND NOT niosII_system_burst_20_upstream_non_bursting_master_requests));
  --niosII_system_burst_20_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_20_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_20_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_20_upstream_arb_share_counter <= niosII_system_burst_20_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_20_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_20_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_20_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_20_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_20_upstream AND NOT niosII_system_burst_20_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_20_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_20_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_20/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_20_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_20_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_20_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_20_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_20/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_20_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_20_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_20_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_20_upstream <= internal_cpu_data_master_requests_niosII_system_burst_20_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_20_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_20_upstream_move_on_to_next_transaction <= niosII_system_burst_20_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_20_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_20_upstream, which is an e_mux
  niosII_system_burst_20_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_20_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --burstcount_fifo_for_niosII_system_burst_20_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_20_upstream : burstcount_fifo_for_niosII_system_burst_20_upstream_module
    port map(
      data_out => niosII_system_burst_20_upstream_transaction_burst_count,
      empty => niosII_system_burst_20_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input78,
      clk => clk,
      data_in => niosII_system_burst_20_upstream_selected_burstcount,
      read => niosII_system_burst_20_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input79,
      write => module_input80
    );

  module_input78 <= std_logic'('0');
  module_input79 <= std_logic'('0');
  module_input80 <= ((in_a_read_cycle AND NOT niosII_system_burst_20_upstream_waits_for_read) AND niosII_system_burst_20_upstream_load_fifo) AND NOT ((niosII_system_burst_20_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_20_upstream_burstcount_fifo_empty));

  --niosII_system_burst_20_upstream current burst minus one, which is an e_assign
  niosII_system_burst_20_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_20_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --what to load in current_burst, for niosII_system_burst_20_upstream, which is an e_mux
  niosII_system_burst_20_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_20_upstream_waits_for_read)) AND NOT niosII_system_burst_20_upstream_load_fifo))) = '1'), (niosII_system_burst_20_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_20_upstream_waits_for_read) AND niosII_system_burst_20_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_20_upstream_burstcount_fifo_empty))) = '1'), (niosII_system_burst_20_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'((niosII_system_burst_20_upstream_this_cycle_is_the_last_burst)) = '1'), (niosII_system_burst_20_upstream_transaction_burst_count & A_ToStdLogicVector(std_logic'('0'))), (std_logic_vector'("0") & (niosII_system_burst_20_upstream_current_burst_minus_one))))), 5);
  --the current burst count for niosII_system_burst_20_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_20_upstream_current_burst <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_20_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_20_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_20_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_20_upstream_current_burst <= niosII_system_burst_20_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_20_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_20_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_20_upstream_waits_for_read)) AND niosII_system_burst_20_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_20_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_20_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_20_upstream_waits_for_read)) AND NOT niosII_system_burst_20_upstream_load_fifo) OR niosII_system_burst_20_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_20_upstream_load_fifo <= p0_niosII_system_burst_20_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_20_upstream, which is an e_assign
  niosII_system_burst_20_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_20_upstream_current_burst_minus_one)) AND niosII_system_burst_20_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_20_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_20_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_20_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_20_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_20_upstream,
      full => open,
      clear_fifo => module_input81,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_20_upstream,
      read => niosII_system_burst_20_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input82,
      write => module_input83
    );

  module_input81 <= std_logic'('0');
  module_input82 <= std_logic'('0');
  module_input83 <= in_a_read_cycle AND NOT niosII_system_burst_20_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_20_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_20_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_20_upstream <= niosII_system_burst_20_upstream_readdatavalid_from_sa;
  --niosII_system_burst_20_upstream_writedata mux, which is an e_mux
  niosII_system_burst_20_upstream_writedata <= cpu_data_master_dbs_write_16;
  --byteaddress mux for niosII_system_burst_20/upstream, which is an e_mux
  niosII_system_burst_20_upstream_byteaddress <= cpu_data_master_address_to_slave (19 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_20_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_20_upstream;
  --cpu/data_master saved-grant niosII_system_burst_20/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_20_upstream <= internal_cpu_data_master_requests_niosII_system_burst_20_upstream;
  --allow new arb cycle for niosII_system_burst_20/upstream, which is an e_assign
  niosII_system_burst_20_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_20_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_20_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_20_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_20_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_20_upstream_begins_xfer) = '1'), niosII_system_burst_20_upstream_unreg_firsttransfer, niosII_system_burst_20_upstream_reg_firsttransfer);
  --niosII_system_burst_20_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_20_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_20_upstream_slavearbiterlockenable AND niosII_system_burst_20_upstream_any_continuerequest));
  --niosII_system_burst_20_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_20_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_20_upstream_begins_xfer) = '1' then 
        niosII_system_burst_20_upstream_reg_firsttransfer <= niosII_system_burst_20_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_20_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_20_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_20_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_20_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_20_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_20_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_20_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_20_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_20_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_20_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_20_upstream_begins_xfer) = '1' then 
        niosII_system_burst_20_upstream_bbt_burstcounter <= niosII_system_burst_20_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_20_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_20_upstream_beginbursttransfer_internal <= niosII_system_burst_20_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_20_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_20_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_20_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_20_upstream AND cpu_data_master_read;
  --niosII_system_burst_20_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_20_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_20_upstream AND cpu_data_master_write;
  --niosII_system_burst_20_upstream_address mux, which is an e_mux
  niosII_system_burst_20_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(cpu_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 19);
  --d1_niosII_system_burst_20_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_20_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_20_upstream_end_xfer <= niosII_system_burst_20_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_20_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_20_upstream_waits_for_read <= niosII_system_burst_20_upstream_in_a_read_cycle AND internal_niosII_system_burst_20_upstream_waitrequest_from_sa;
  --niosII_system_burst_20_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_20_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_20_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_20_upstream_in_a_read_cycle;
  --niosII_system_burst_20_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_20_upstream_waits_for_write <= niosII_system_burst_20_upstream_in_a_write_cycle AND internal_niosII_system_burst_20_upstream_waitrequest_from_sa;
  --niosII_system_burst_20_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_20_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_20_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_20_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_20_upstream_counter <= std_logic'('0');
  --niosII_system_burst_20_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_20_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_20_upstream)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_byteenable_niosII_system_burst_20_upstream)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  (cpu_data_master_byteenable_niosII_system_burst_20_upstream_segment_1(1), cpu_data_master_byteenable_niosII_system_burst_20_upstream_segment_1(0), cpu_data_master_byteenable_niosII_system_burst_20_upstream_segment_0(1), cpu_data_master_byteenable_niosII_system_burst_20_upstream_segment_0(0)) <= cpu_data_master_byteenable;
  internal_cpu_data_master_byteenable_niosII_system_burst_20_upstream <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), cpu_data_master_byteenable_niosII_system_burst_20_upstream_segment_0, cpu_data_master_byteenable_niosII_system_burst_20_upstream_segment_1);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_20_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_20_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_20_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_20_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_byteenable_niosII_system_burst_20_upstream <= internal_cpu_data_master_byteenable_niosII_system_burst_20_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_20_upstream <= internal_cpu_data_master_granted_niosII_system_burst_20_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_20_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_20_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_20_upstream <= internal_cpu_data_master_requests_niosII_system_burst_20_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_20_upstream_burstcount <= internal_niosII_system_burst_20_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_20_upstream_read <= internal_niosII_system_burst_20_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_20_upstream_waitrequest_from_sa <= internal_niosII_system_burst_20_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_20_upstream_write <= internal_niosII_system_burst_20_upstream_write;
--synthesis translate_off
    --niosII_system_burst_20/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line122 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_20_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line122, now);
          write(write_line122, string'(": "));
          write(write_line122, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_20/upstream"));
          write(output, write_line122.all);
          deallocate (write_line122);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_20_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_tsb_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal incoming_sram_IF_0_tsb_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_address : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_20_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_granted_sram_IF_0_tsb : IN STD_LOGIC;
                 signal niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb : IN STD_LOGIC;
                 signal niosII_system_burst_20_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb : IN STD_LOGIC;
                 signal niosII_system_burst_20_downstream_requests_sram_IF_0_tsb : IN STD_LOGIC;
                 signal niosII_system_burst_20_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_20_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_20_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_20_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_20_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_20_downstream_arbitrator;


architecture europa of niosII_system_burst_20_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_20_downstream_address_to_slave :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal internal_niosII_system_burst_20_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_niosII_system_burst_20_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_20_downstream_address_last_time :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_20_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_20_downstream_is_granted_some_slave :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_niosII_system_burst_20_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pre_flush_niosII_system_burst_20_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb OR NOT niosII_system_burst_20_downstream_requests_sram_IF_0_tsb)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_20_downstream_granted_sram_IF_0_tsb OR NOT niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb OR NOT niosII_system_burst_20_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_tsb_avalon_slave_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_20_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb OR NOT niosII_system_burst_20_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_20_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_20_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_20_downstream_address_to_slave <= niosII_system_burst_20_downstream_address;
  --niosII_system_burst_20_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_20_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_20_downstream_read_but_no_slave_selected <= (niosII_system_burst_20_downstream_read AND niosII_system_burst_20_downstream_run) AND NOT niosII_system_burst_20_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  niosII_system_burst_20_downstream_is_granted_some_slave <= niosII_system_burst_20_downstream_granted_sram_IF_0_tsb;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_20_downstream_readdatavalid <= niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb;
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_20_downstream_readdatavalid <= niosII_system_burst_20_downstream_read_but_no_slave_selected OR pre_flush_niosII_system_burst_20_downstream_readdatavalid;
  --niosII_system_burst_20/downstream readdata mux, which is an e_mux
  niosII_system_burst_20_downstream_readdata <= incoming_sram_IF_0_tsb_data;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_20_downstream_waitrequest <= NOT niosII_system_burst_20_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_niosII_system_burst_20_downstream_latency_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      internal_niosII_system_burst_20_downstream_latency_counter <= p1_niosII_system_burst_20_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_niosII_system_burst_20_downstream_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((niosII_system_burst_20_downstream_run AND niosII_system_burst_20_downstream_read))) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_niosII_system_burst_20_downstream_latency_counter)) /= std_logic_vector'("00")), ((std_logic_vector'("0000000000000000000000000000000") & (internal_niosII_system_burst_20_downstream_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (A_REP(niosII_system_burst_20_downstream_requests_sram_IF_0_tsb, 2))) AND std_logic_vector'("00000000000000000000000000000010")), 2);
  --niosII_system_burst_20_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_20_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_20_downstream_address_to_slave <= internal_niosII_system_burst_20_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_20_downstream_latency_counter <= internal_niosII_system_burst_20_downstream_latency_counter;
  --vhdl renameroo for output signals
  niosII_system_burst_20_downstream_waitrequest <= internal_niosII_system_burst_20_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_20_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_20_downstream_address_last_time <= std_logic_vector'("0000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_20_downstream_address_last_time <= niosII_system_burst_20_downstream_address;
      end if;

    end process;

    --niosII_system_burst_20/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_20_downstream_waitrequest AND ((niosII_system_burst_20_downstream_read OR niosII_system_burst_20_downstream_write));
      end if;

    end process;

    --niosII_system_burst_20_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line123 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_20_downstream_address /= niosII_system_burst_20_downstream_address_last_time))))) = '1' then 
          write(write_line123, now);
          write(write_line123, string'(": "));
          write(write_line123, string'("niosII_system_burst_20_downstream_address did not heed wait!!!"));
          write(output, write_line123.all);
          deallocate (write_line123);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_20_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_20_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_20_downstream_burstcount_last_time <= niosII_system_burst_20_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_20_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line124 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_20_downstream_burstcount) /= std_logic'(niosII_system_burst_20_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line124, now);
          write(write_line124, string'(": "));
          write(write_line124, string'("niosII_system_burst_20_downstream_burstcount did not heed wait!!!"));
          write(output, write_line124.all);
          deallocate (write_line124);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_20_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_20_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_20_downstream_byteenable_last_time <= niosII_system_burst_20_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_20_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line125 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_20_downstream_byteenable /= niosII_system_burst_20_downstream_byteenable_last_time))))) = '1' then 
          write(write_line125, now);
          write(write_line125, string'(": "));
          write(write_line125, string'("niosII_system_burst_20_downstream_byteenable did not heed wait!!!"));
          write(output, write_line125.all);
          deallocate (write_line125);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_20_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_20_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_20_downstream_read_last_time <= niosII_system_burst_20_downstream_read;
      end if;

    end process;

    --niosII_system_burst_20_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line126 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_20_downstream_read) /= std_logic'(niosII_system_burst_20_downstream_read_last_time)))))) = '1' then 
          write(write_line126, now);
          write(write_line126, string'(": "));
          write(write_line126, string'("niosII_system_burst_20_downstream_read did not heed wait!!!"));
          write(output, write_line126.all);
          deallocate (write_line126);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_20_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_20_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_20_downstream_write_last_time <= niosII_system_burst_20_downstream_write;
      end if;

    end process;

    --niosII_system_burst_20_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line127 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_20_downstream_write) /= std_logic'(niosII_system_burst_20_downstream_write_last_time)))))) = '1' then 
          write(write_line127, now);
          write(write_line127, string'(": "));
          write(write_line127, string'("niosII_system_burst_20_downstream_write did not heed wait!!!"));
          write(output, write_line127.all);
          deallocate (write_line127);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_20_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_20_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_20_downstream_writedata_last_time <= niosII_system_burst_20_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_20_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line128 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_20_downstream_writedata /= niosII_system_burst_20_downstream_writedata_last_time)))) AND niosII_system_burst_20_downstream_write)) = '1' then 
          write(write_line128, now);
          write(write_line128, string'(": "));
          write(write_line128, string'("niosII_system_burst_20_downstream_writedata did not heed wait!!!"));
          write(output, write_line128.all);
          deallocate (write_line128);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_21_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_21_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_21_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_21_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_21_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_21_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_21_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_21_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_21_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_21_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_21_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_21_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_21_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_21_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_21_upstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_21_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_21_upstream_byteaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal niosII_system_burst_21_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_21_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_21_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_21_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_21_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_21_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_21_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity niosII_system_burst_21_upstream_arbitrator;


architecture europa of niosII_system_burst_21_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_21_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_21_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_21_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_21_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_21_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_21_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_21_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_21_upstream_write :  STD_LOGIC;
                signal module_input84 :  STD_LOGIC;
                signal module_input85 :  STD_LOGIC;
                signal module_input86 :  STD_LOGIC;
                signal module_input87 :  STD_LOGIC;
                signal module_input88 :  STD_LOGIC;
                signal module_input89 :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_21_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_21_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_21_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_21_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_21_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_21_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_21_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_21_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_21_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_21_upstream);
  --assign niosII_system_burst_21_upstream_readdatavalid_from_sa = niosII_system_burst_21_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_21_upstream_readdatavalid_from_sa <= niosII_system_burst_21_upstream_readdatavalid;
  --assign niosII_system_burst_21_upstream_readdata_from_sa = niosII_system_burst_21_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_21_upstream_readdata_from_sa <= niosII_system_burst_21_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_21_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1100100001001000010110000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_21_upstream_waitrequest_from_sa = niosII_system_burst_21_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_21_upstream_waitrequest_from_sa <= niosII_system_burst_21_upstream_waitrequest;
  --niosII_system_burst_21_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_21_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_21_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_21_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_21_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_21_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_21_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_21_upstream;
  --niosII_system_burst_21_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_21_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_21_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_21_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_21_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_21_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_21_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_21_upstream_allgrants <= niosII_system_burst_21_upstream_grant_vector;
  --niosII_system_burst_21_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_21_upstream_end_xfer <= NOT ((niosII_system_burst_21_upstream_waits_for_read OR niosII_system_burst_21_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_21_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_21_upstream <= niosII_system_burst_21_upstream_end_xfer AND (((NOT niosII_system_burst_21_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_21_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_21_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_21_upstream AND niosII_system_burst_21_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_21_upstream AND NOT niosII_system_burst_21_upstream_non_bursting_master_requests));
  --niosII_system_burst_21_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_21_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_21_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_21_upstream_arb_share_counter <= niosII_system_burst_21_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_21_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_21_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_21_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_21_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_21_upstream AND NOT niosII_system_burst_21_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_21_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_21_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_21/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_21_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_21_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_21_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_21_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_21/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_21_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_21_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_21_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_21_upstream <= internal_cpu_data_master_requests_niosII_system_burst_21_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_21_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_21_upstream_move_on_to_next_transaction <= niosII_system_burst_21_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_21_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_21_upstream, which is an e_mux
  niosII_system_burst_21_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_21_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_21_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_21_upstream : burstcount_fifo_for_niosII_system_burst_21_upstream_module
    port map(
      data_out => niosII_system_burst_21_upstream_transaction_burst_count,
      empty => niosII_system_burst_21_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input84,
      clk => clk,
      data_in => niosII_system_burst_21_upstream_selected_burstcount,
      read => niosII_system_burst_21_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input85,
      write => module_input86
    );

  module_input84 <= std_logic'('0');
  module_input85 <= std_logic'('0');
  module_input86 <= ((in_a_read_cycle AND NOT niosII_system_burst_21_upstream_waits_for_read) AND niosII_system_burst_21_upstream_load_fifo) AND NOT ((niosII_system_burst_21_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_21_upstream_burstcount_fifo_empty));

  --niosII_system_burst_21_upstream current burst minus one, which is an e_assign
  niosII_system_burst_21_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_21_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_21_upstream, which is an e_mux
  niosII_system_burst_21_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_21_upstream_waits_for_read)) AND NOT niosII_system_burst_21_upstream_load_fifo))) = '1'), niosII_system_burst_21_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_21_upstream_waits_for_read) AND niosII_system_burst_21_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_21_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_21_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_21_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_21_upstream_transaction_burst_count, niosII_system_burst_21_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_21_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_21_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_21_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_21_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_21_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_21_upstream_current_burst <= niosII_system_burst_21_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_21_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_21_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_21_upstream_waits_for_read)) AND niosII_system_burst_21_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_21_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_21_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_21_upstream_waits_for_read)) AND NOT niosII_system_burst_21_upstream_load_fifo) OR niosII_system_burst_21_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_21_upstream_load_fifo <= p0_niosII_system_burst_21_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_21_upstream, which is an e_assign
  niosII_system_burst_21_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_21_upstream_current_burst_minus_one)) AND niosII_system_burst_21_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_21_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_21_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_21_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_21_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_21_upstream,
      full => open,
      clear_fifo => module_input87,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_21_upstream,
      read => niosII_system_burst_21_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input88,
      write => module_input89
    );

  module_input87 <= std_logic'('0');
  module_input88 <= std_logic'('0');
  module_input89 <= in_a_read_cycle AND NOT niosII_system_burst_21_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_21_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_21_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_21_upstream <= niosII_system_burst_21_upstream_readdatavalid_from_sa;
  --niosII_system_burst_21_upstream_writedata mux, which is an e_mux
  niosII_system_burst_21_upstream_writedata <= cpu_data_master_writedata;
  --byteaddress mux for niosII_system_burst_21/upstream, which is an e_mux
  niosII_system_burst_21_upstream_byteaddress <= cpu_data_master_address_to_slave (5 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_21_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_21_upstream;
  --cpu/data_master saved-grant niosII_system_burst_21/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_21_upstream <= internal_cpu_data_master_requests_niosII_system_burst_21_upstream;
  --allow new arb cycle for niosII_system_burst_21/upstream, which is an e_assign
  niosII_system_burst_21_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_21_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_21_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_21_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_21_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_21_upstream_begins_xfer) = '1'), niosII_system_burst_21_upstream_unreg_firsttransfer, niosII_system_burst_21_upstream_reg_firsttransfer);
  --niosII_system_burst_21_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_21_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_21_upstream_slavearbiterlockenable AND niosII_system_burst_21_upstream_any_continuerequest));
  --niosII_system_burst_21_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_21_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_21_upstream_begins_xfer) = '1' then 
        niosII_system_burst_21_upstream_reg_firsttransfer <= niosII_system_burst_21_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_21_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_21_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_21_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_21_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_21_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_21_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_21_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_21_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_21_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_21_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_21_upstream_begins_xfer) = '1' then 
        niosII_system_burst_21_upstream_bbt_burstcounter <= niosII_system_burst_21_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_21_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_21_upstream_beginbursttransfer_internal <= niosII_system_burst_21_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_21_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_21_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_21_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_21_upstream AND cpu_data_master_read;
  --niosII_system_burst_21_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_21_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_21_upstream AND cpu_data_master_write;
  --niosII_system_burst_21_upstream_address mux, which is an e_mux
  niosII_system_burst_21_upstream_address <= cpu_data_master_address_to_slave (3 DOWNTO 0);
  --d1_niosII_system_burst_21_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_21_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_21_upstream_end_xfer <= niosII_system_burst_21_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_21_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_21_upstream_waits_for_read <= niosII_system_burst_21_upstream_in_a_read_cycle AND internal_niosII_system_burst_21_upstream_waitrequest_from_sa;
  --niosII_system_burst_21_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_21_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_21_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_21_upstream_in_a_read_cycle;
  --niosII_system_burst_21_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_21_upstream_waits_for_write <= niosII_system_burst_21_upstream_in_a_write_cycle AND internal_niosII_system_burst_21_upstream_waitrequest_from_sa;
  --niosII_system_burst_21_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_21_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_21_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_21_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_21_upstream_counter <= std_logic'('0');
  --niosII_system_burst_21_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_21_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_21_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_21_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_21_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_21_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_21_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_21_upstream <= internal_cpu_data_master_granted_niosII_system_burst_21_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_21_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_21_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_21_upstream <= internal_cpu_data_master_requests_niosII_system_burst_21_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_21_upstream_burstcount <= internal_niosII_system_burst_21_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_21_upstream_read <= internal_niosII_system_burst_21_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_21_upstream_waitrequest_from_sa <= internal_niosII_system_burst_21_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_21_upstream_write <= internal_niosII_system_burst_21_upstream_write;
--synthesis translate_off
    --niosII_system_burst_21/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line129 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_21_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line129, now);
          write(write_line129, string'(": "));
          write(write_line129, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_21/upstream"));
          write(output, write_line129.all);
          deallocate (write_line129);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_21_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_niosII_system_clock_0_in_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_21_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_21_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_21_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_21_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_21_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_21_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_21_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_21_downstream_arbitrator;


architecture europa of niosII_system_burst_21_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_21_downstream_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_21_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_flush_niosII_system_burst_21_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in OR NOT niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in OR NOT ((niosII_system_burst_21_downstream_read OR niosII_system_burst_21_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_21_downstream_read OR niosII_system_burst_21_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in OR NOT ((niosII_system_burst_21_downstream_read OR niosII_system_burst_21_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_21_downstream_read OR niosII_system_burst_21_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_21_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_21_downstream_address_to_slave <= niosII_system_burst_21_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_21_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_21_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_21_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in)))));
  --niosII_system_burst_21/downstream readdata mux, which is an e_mux
  niosII_system_burst_21_downstream_readdata <= niosII_system_clock_0_in_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_21_downstream_waitrequest <= NOT niosII_system_burst_21_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_21_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_21_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_21_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_21_downstream_address_to_slave <= internal_niosII_system_burst_21_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_21_downstream_waitrequest <= internal_niosII_system_burst_21_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_21_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_21_downstream_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_21_downstream_address_last_time <= niosII_system_burst_21_downstream_address;
      end if;

    end process;

    --niosII_system_burst_21/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_21_downstream_waitrequest AND ((niosII_system_burst_21_downstream_read OR niosII_system_burst_21_downstream_write));
      end if;

    end process;

    --niosII_system_burst_21_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line130 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_21_downstream_address /= niosII_system_burst_21_downstream_address_last_time))))) = '1' then 
          write(write_line130, now);
          write(write_line130, string'(": "));
          write(write_line130, string'("niosII_system_burst_21_downstream_address did not heed wait!!!"));
          write(output, write_line130.all);
          deallocate (write_line130);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_21_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_21_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_21_downstream_burstcount_last_time <= niosII_system_burst_21_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_21_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line131 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_21_downstream_burstcount) /= std_logic'(niosII_system_burst_21_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line131, now);
          write(write_line131, string'(": "));
          write(write_line131, string'("niosII_system_burst_21_downstream_burstcount did not heed wait!!!"));
          write(output, write_line131.all);
          deallocate (write_line131);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_21_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_21_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_21_downstream_byteenable_last_time <= niosII_system_burst_21_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_21_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line132 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_21_downstream_byteenable /= niosII_system_burst_21_downstream_byteenable_last_time))))) = '1' then 
          write(write_line132, now);
          write(write_line132, string'(": "));
          write(write_line132, string'("niosII_system_burst_21_downstream_byteenable did not heed wait!!!"));
          write(output, write_line132.all);
          deallocate (write_line132);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_21_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_21_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_21_downstream_read_last_time <= niosII_system_burst_21_downstream_read;
      end if;

    end process;

    --niosII_system_burst_21_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line133 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_21_downstream_read) /= std_logic'(niosII_system_burst_21_downstream_read_last_time)))))) = '1' then 
          write(write_line133, now);
          write(write_line133, string'(": "));
          write(write_line133, string'("niosII_system_burst_21_downstream_read did not heed wait!!!"));
          write(output, write_line133.all);
          deallocate (write_line133);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_21_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_21_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_21_downstream_write_last_time <= niosII_system_burst_21_downstream_write;
      end if;

    end process;

    --niosII_system_burst_21_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line134 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_21_downstream_write) /= std_logic'(niosII_system_burst_21_downstream_write_last_time)))))) = '1' then 
          write(write_line134, now);
          write(write_line134, string'(": "));
          write(write_line134, string'("niosII_system_burst_21_downstream_write did not heed wait!!!"));
          write(output, write_line134.all);
          deallocate (write_line134);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_21_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_21_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_21_downstream_writedata_last_time <= niosII_system_burst_21_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_21_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line135 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_21_downstream_writedata /= niosII_system_burst_21_downstream_writedata_last_time)))) AND niosII_system_burst_21_downstream_write)) = '1' then 
          write(write_line135, now);
          write(write_line135, string'(": "));
          write(write_line135, string'("niosII_system_burst_21_downstream_writedata did not heed wait!!!"));
          write(output, write_line135.all);
          deallocate (write_line135);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_3_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_3_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_3_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("0000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_3_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_3_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_3_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_3_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_3_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_3_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_3_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_3_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_3_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_3_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_3_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_3_upstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal niosII_system_burst_3_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_3_upstream_byteaddress : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_3_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_3_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_3_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_3_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_3_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_3_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_3_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity niosII_system_burst_3_upstream_arbitrator;


architecture europa of niosII_system_burst_3_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_3_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_3_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_3_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_3_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_3_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_3_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_3_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_3_upstream_write :  STD_LOGIC;
                signal module_input90 :  STD_LOGIC;
                signal module_input91 :  STD_LOGIC;
                signal module_input92 :  STD_LOGIC;
                signal module_input93 :  STD_LOGIC;
                signal module_input94 :  STD_LOGIC;
                signal module_input95 :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_3_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_3_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_3_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_3_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_3_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_3_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_3_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_3_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_3_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_3_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_3_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_niosII_system_burst_3_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_3_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_3_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_3_upstream);
  --assign niosII_system_burst_3_upstream_readdatavalid_from_sa = niosII_system_burst_3_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_3_upstream_readdatavalid_from_sa <= niosII_system_burst_3_upstream_readdatavalid;
  --assign niosII_system_burst_3_upstream_readdata_from_sa = niosII_system_burst_3_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_3_upstream_readdata_from_sa <= niosII_system_burst_3_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_3_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 14) & std_logic_vector'("00000000000000")) = std_logic_vector'("1100100000100000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_3_upstream_waitrequest_from_sa = niosII_system_burst_3_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_3_upstream_waitrequest_from_sa <= niosII_system_burst_3_upstream_waitrequest;
  --niosII_system_burst_3_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_3_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_3_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_3_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_3_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_3_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_3_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_3_upstream;
  --niosII_system_burst_3_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_3_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_3_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_3_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_3_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_3_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_3_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_3_upstream_allgrants <= niosII_system_burst_3_upstream_grant_vector;
  --niosII_system_burst_3_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_3_upstream_end_xfer <= NOT ((niosII_system_burst_3_upstream_waits_for_read OR niosII_system_burst_3_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_3_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_3_upstream <= niosII_system_burst_3_upstream_end_xfer AND (((NOT niosII_system_burst_3_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_3_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_3_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_3_upstream AND niosII_system_burst_3_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_3_upstream AND NOT niosII_system_burst_3_upstream_non_bursting_master_requests));
  --niosII_system_burst_3_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_3_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_3_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_3_upstream_arb_share_counter <= niosII_system_burst_3_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_3_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_3_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_3_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_3_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_3_upstream AND NOT niosII_system_burst_3_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_3_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_3_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_3/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_3_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_3_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_3_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_3_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_3/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_3_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_3_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_3_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_3_upstream <= internal_cpu_data_master_requests_niosII_system_burst_3_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_3_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_3_upstream_move_on_to_next_transaction <= niosII_system_burst_3_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_3_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_3_upstream, which is an e_mux
  niosII_system_burst_3_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_3_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_3_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_3_upstream : burstcount_fifo_for_niosII_system_burst_3_upstream_module
    port map(
      data_out => niosII_system_burst_3_upstream_transaction_burst_count,
      empty => niosII_system_burst_3_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input90,
      clk => clk,
      data_in => niosII_system_burst_3_upstream_selected_burstcount,
      read => niosII_system_burst_3_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input91,
      write => module_input92
    );

  module_input90 <= std_logic'('0');
  module_input91 <= std_logic'('0');
  module_input92 <= ((in_a_read_cycle AND NOT niosII_system_burst_3_upstream_waits_for_read) AND niosII_system_burst_3_upstream_load_fifo) AND NOT ((niosII_system_burst_3_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_3_upstream_burstcount_fifo_empty));

  --niosII_system_burst_3_upstream current burst minus one, which is an e_assign
  niosII_system_burst_3_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_3_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_3_upstream, which is an e_mux
  niosII_system_burst_3_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_3_upstream_waits_for_read)) AND NOT niosII_system_burst_3_upstream_load_fifo))) = '1'), niosII_system_burst_3_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_3_upstream_waits_for_read) AND niosII_system_burst_3_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_3_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_3_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_3_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_3_upstream_transaction_burst_count, niosII_system_burst_3_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_3_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_3_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_3_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_3_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_3_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_3_upstream_current_burst <= niosII_system_burst_3_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_3_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_3_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_3_upstream_waits_for_read)) AND niosII_system_burst_3_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_3_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_3_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_3_upstream_waits_for_read)) AND NOT niosII_system_burst_3_upstream_load_fifo) OR niosII_system_burst_3_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_3_upstream_load_fifo <= p0_niosII_system_burst_3_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_3_upstream, which is an e_assign
  niosII_system_burst_3_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_3_upstream_current_burst_minus_one)) AND niosII_system_burst_3_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_3_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_3_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_3_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_3_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_3_upstream,
      full => open,
      clear_fifo => module_input93,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_3_upstream,
      read => niosII_system_burst_3_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input94,
      write => module_input95
    );

  module_input93 <= std_logic'('0');
  module_input94 <= std_logic'('0');
  module_input95 <= in_a_read_cycle AND NOT niosII_system_burst_3_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_3_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_3_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_3_upstream <= niosII_system_burst_3_upstream_readdatavalid_from_sa;
  --niosII_system_burst_3_upstream_writedata mux, which is an e_mux
  niosII_system_burst_3_upstream_writedata <= cpu_data_master_writedata;
  --byteaddress mux for niosII_system_burst_3/upstream, which is an e_mux
  niosII_system_burst_3_upstream_byteaddress <= cpu_data_master_address_to_slave (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_3_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_3_upstream;
  --cpu/data_master saved-grant niosII_system_burst_3/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_3_upstream <= internal_cpu_data_master_requests_niosII_system_burst_3_upstream;
  --allow new arb cycle for niosII_system_burst_3/upstream, which is an e_assign
  niosII_system_burst_3_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_3_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_3_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_3_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_3_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_3_upstream_begins_xfer) = '1'), niosII_system_burst_3_upstream_unreg_firsttransfer, niosII_system_burst_3_upstream_reg_firsttransfer);
  --niosII_system_burst_3_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_3_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_3_upstream_slavearbiterlockenable AND niosII_system_burst_3_upstream_any_continuerequest));
  --niosII_system_burst_3_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_3_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_3_upstream_begins_xfer) = '1' then 
        niosII_system_burst_3_upstream_reg_firsttransfer <= niosII_system_burst_3_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_3_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_3_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_3_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_3_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_3_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_3_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_3_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_3_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_3_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_3_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_3_upstream_begins_xfer) = '1' then 
        niosII_system_burst_3_upstream_bbt_burstcounter <= niosII_system_burst_3_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_3_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_3_upstream_beginbursttransfer_internal <= niosII_system_burst_3_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_3_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_3_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_3_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_3_upstream AND cpu_data_master_read;
  --niosII_system_burst_3_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_3_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_3_upstream AND cpu_data_master_write;
  --niosII_system_burst_3_upstream_address mux, which is an e_mux
  niosII_system_burst_3_upstream_address <= cpu_data_master_address_to_slave (13 DOWNTO 0);
  --d1_niosII_system_burst_3_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_3_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_3_upstream_end_xfer <= niosII_system_burst_3_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_3_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_3_upstream_waits_for_read <= niosII_system_burst_3_upstream_in_a_read_cycle AND internal_niosII_system_burst_3_upstream_waitrequest_from_sa;
  --niosII_system_burst_3_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_3_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_3_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_3_upstream_in_a_read_cycle;
  --niosII_system_burst_3_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_3_upstream_waits_for_write <= niosII_system_burst_3_upstream_in_a_write_cycle AND internal_niosII_system_burst_3_upstream_waitrequest_from_sa;
  --niosII_system_burst_3_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_3_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_3_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_3_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_3_upstream_counter <= std_logic'('0');
  --niosII_system_burst_3_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_3_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_3_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_3_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_3_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_3_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_3_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_3_upstream <= internal_cpu_data_master_granted_niosII_system_burst_3_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_3_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_3_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_3_upstream <= internal_cpu_data_master_requests_niosII_system_burst_3_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_3_upstream_burstcount <= internal_niosII_system_burst_3_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_3_upstream_read <= internal_niosII_system_burst_3_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_3_upstream_waitrequest_from_sa <= internal_niosII_system_burst_3_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_3_upstream_write <= internal_niosII_system_burst_3_upstream_write;
--synthesis translate_off
    --niosII_system_burst_3/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line136 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_3_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line136, now);
          write(write_line136, string'(": "));
          write(write_line136, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_3/upstream"));
          write(output, write_line136.all);
          deallocate (write_line136);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_3_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_memory_s1_end_xfer : IN STD_LOGIC;
                 signal memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_3_downstream_address : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal niosII_system_burst_3_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_3_downstream_granted_memory_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_qualified_request_memory_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_read_data_valid_memory_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_requests_memory_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_3_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal niosII_system_burst_3_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_3_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_3_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_3_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_3_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_3_downstream_arbitrator;


architecture europa of niosII_system_burst_3_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_3_downstream_address_to_slave :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal internal_niosII_system_burst_3_downstream_latency_counter :  STD_LOGIC;
                signal internal_niosII_system_burst_3_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_address_last_time :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_3_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_3_downstream_is_granted_some_slave :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_niosII_system_burst_3_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_niosII_system_burst_3_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_3_downstream_qualified_request_memory_s1 OR NOT niosII_system_burst_3_downstream_requests_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_3_downstream_granted_memory_s1 OR NOT niosII_system_burst_3_downstream_qualified_request_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_3_downstream_qualified_request_memory_s1 OR NOT ((niosII_system_burst_3_downstream_read OR niosII_system_burst_3_downstream_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_3_downstream_read OR niosII_system_burst_3_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_3_downstream_qualified_request_memory_s1 OR NOT ((niosII_system_burst_3_downstream_read OR niosII_system_burst_3_downstream_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_3_downstream_read OR niosII_system_burst_3_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_3_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_3_downstream_address_to_slave <= niosII_system_burst_3_downstream_address;
  --niosII_system_burst_3_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_3_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      niosII_system_burst_3_downstream_read_but_no_slave_selected <= (niosII_system_burst_3_downstream_read AND niosII_system_burst_3_downstream_run) AND NOT niosII_system_burst_3_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  niosII_system_burst_3_downstream_is_granted_some_slave <= niosII_system_burst_3_downstream_granted_memory_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_3_downstream_readdatavalid <= niosII_system_burst_3_downstream_read_data_valid_memory_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_3_downstream_readdatavalid <= niosII_system_burst_3_downstream_read_but_no_slave_selected OR pre_flush_niosII_system_burst_3_downstream_readdatavalid;
  --niosII_system_burst_3/downstream readdata mux, which is an e_mux
  niosII_system_burst_3_downstream_readdata <= memory_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_3_downstream_waitrequest <= NOT niosII_system_burst_3_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_niosII_system_burst_3_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_niosII_system_burst_3_downstream_latency_counter <= p1_niosII_system_burst_3_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_niosII_system_burst_3_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((niosII_system_burst_3_downstream_run AND niosII_system_burst_3_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_3_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_3_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_3_downstream_requests_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --niosII_system_burst_3_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_3_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_3_downstream_address_to_slave <= internal_niosII_system_burst_3_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_3_downstream_latency_counter <= internal_niosII_system_burst_3_downstream_latency_counter;
  --vhdl renameroo for output signals
  niosII_system_burst_3_downstream_waitrequest <= internal_niosII_system_burst_3_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_3_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_3_downstream_address_last_time <= std_logic_vector'("00000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_3_downstream_address_last_time <= niosII_system_burst_3_downstream_address;
      end if;

    end process;

    --niosII_system_burst_3/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_3_downstream_waitrequest AND ((niosII_system_burst_3_downstream_read OR niosII_system_burst_3_downstream_write));
      end if;

    end process;

    --niosII_system_burst_3_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line137 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_3_downstream_address /= niosII_system_burst_3_downstream_address_last_time))))) = '1' then 
          write(write_line137, now);
          write(write_line137, string'(": "));
          write(write_line137, string'("niosII_system_burst_3_downstream_address did not heed wait!!!"));
          write(output, write_line137.all);
          deallocate (write_line137);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_3_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_3_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_3_downstream_burstcount_last_time <= niosII_system_burst_3_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_3_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line138 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_3_downstream_burstcount) /= std_logic'(niosII_system_burst_3_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line138, now);
          write(write_line138, string'(": "));
          write(write_line138, string'("niosII_system_burst_3_downstream_burstcount did not heed wait!!!"));
          write(output, write_line138.all);
          deallocate (write_line138);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_3_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_3_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_3_downstream_byteenable_last_time <= niosII_system_burst_3_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_3_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line139 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_3_downstream_byteenable /= niosII_system_burst_3_downstream_byteenable_last_time))))) = '1' then 
          write(write_line139, now);
          write(write_line139, string'(": "));
          write(write_line139, string'("niosII_system_burst_3_downstream_byteenable did not heed wait!!!"));
          write(output, write_line139.all);
          deallocate (write_line139);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_3_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_3_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_3_downstream_read_last_time <= niosII_system_burst_3_downstream_read;
      end if;

    end process;

    --niosII_system_burst_3_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line140 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_3_downstream_read) /= std_logic'(niosII_system_burst_3_downstream_read_last_time)))))) = '1' then 
          write(write_line140, now);
          write(write_line140, string'(": "));
          write(write_line140, string'("niosII_system_burst_3_downstream_read did not heed wait!!!"));
          write(output, write_line140.all);
          deallocate (write_line140);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_3_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_3_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_3_downstream_write_last_time <= niosII_system_burst_3_downstream_write;
      end if;

    end process;

    --niosII_system_burst_3_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line141 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_3_downstream_write) /= std_logic'(niosII_system_burst_3_downstream_write_last_time)))))) = '1' then 
          write(write_line141, now);
          write(write_line141, string'(": "));
          write(write_line141, string'("niosII_system_burst_3_downstream_write did not heed wait!!!"));
          write(output, write_line141.all);
          deallocate (write_line141);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_3_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_3_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_3_downstream_writedata_last_time <= niosII_system_burst_3_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_3_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line142 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_3_downstream_writedata /= niosII_system_burst_3_downstream_writedata_last_time)))) AND niosII_system_burst_3_downstream_write)) = '1' then 
          write(write_line142, now);
          write(write_line142, string'(": "));
          write(write_line142, string'("niosII_system_burst_3_downstream_writedata did not heed wait!!!"));
          write(output, write_line142.all);
          deallocate (write_line142);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_4_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_4_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_4_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_4_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_4_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_4_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_4_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_4_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_4_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_4_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_4_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_4_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_4_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_4_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_4_upstream_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_4_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_4_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_4_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_4_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_4_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_4_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_4_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_4_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_4_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity niosII_system_burst_4_upstream_arbitrator;


architecture europa of niosII_system_burst_4_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_4_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_4_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_4_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_4_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_4_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_4_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_4_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_4_upstream_write :  STD_LOGIC;
                signal module_input100 :  STD_LOGIC;
                signal module_input101 :  STD_LOGIC;
                signal module_input96 :  STD_LOGIC;
                signal module_input97 :  STD_LOGIC;
                signal module_input98 :  STD_LOGIC;
                signal module_input99 :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_4_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_4_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_4_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_4_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_4_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_4_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_4_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_4_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_4_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_4_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_4_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_4_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_4_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_4_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_4_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_4_upstream);
  --assign niosII_system_burst_4_upstream_readdatavalid_from_sa = niosII_system_burst_4_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_4_upstream_readdatavalid_from_sa <= niosII_system_burst_4_upstream_readdatavalid;
  --assign niosII_system_burst_4_upstream_readdata_from_sa = niosII_system_burst_4_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_4_upstream_readdata_from_sa <= niosII_system_burst_4_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_4_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("1100100001001000011010000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_4_upstream_waitrequest_from_sa = niosII_system_burst_4_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_4_upstream_waitrequest_from_sa <= niosII_system_burst_4_upstream_waitrequest;
  --niosII_system_burst_4_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_4_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_4_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_4_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_4_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_4_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_4_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_4_upstream;
  --niosII_system_burst_4_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_4_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_4_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_4_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_4_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_4_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_4_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_4_upstream_allgrants <= niosII_system_burst_4_upstream_grant_vector;
  --niosII_system_burst_4_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_4_upstream_end_xfer <= NOT ((niosII_system_burst_4_upstream_waits_for_read OR niosII_system_burst_4_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_4_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_4_upstream <= niosII_system_burst_4_upstream_end_xfer AND (((NOT niosII_system_burst_4_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_4_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_4_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_4_upstream AND niosII_system_burst_4_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_4_upstream AND NOT niosII_system_burst_4_upstream_non_bursting_master_requests));
  --niosII_system_burst_4_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_4_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_4_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_4_upstream_arb_share_counter <= niosII_system_burst_4_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_4_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_4_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_4_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_4_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_4_upstream AND NOT niosII_system_burst_4_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_4_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_4_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_4/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_4_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_4_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_4_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_4_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_4/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_4_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_4_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_4_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_4_upstream <= internal_cpu_data_master_requests_niosII_system_burst_4_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_4_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_4_upstream_move_on_to_next_transaction <= niosII_system_burst_4_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_4_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_4_upstream, which is an e_mux
  niosII_system_burst_4_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_4_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_4_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_4_upstream : burstcount_fifo_for_niosII_system_burst_4_upstream_module
    port map(
      data_out => niosII_system_burst_4_upstream_transaction_burst_count,
      empty => niosII_system_burst_4_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input96,
      clk => clk,
      data_in => niosII_system_burst_4_upstream_selected_burstcount,
      read => niosII_system_burst_4_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input97,
      write => module_input98
    );

  module_input96 <= std_logic'('0');
  module_input97 <= std_logic'('0');
  module_input98 <= ((in_a_read_cycle AND NOT niosII_system_burst_4_upstream_waits_for_read) AND niosII_system_burst_4_upstream_load_fifo) AND NOT ((niosII_system_burst_4_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_4_upstream_burstcount_fifo_empty));

  --niosII_system_burst_4_upstream current burst minus one, which is an e_assign
  niosII_system_burst_4_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_4_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_4_upstream, which is an e_mux
  niosII_system_burst_4_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_4_upstream_waits_for_read)) AND NOT niosII_system_burst_4_upstream_load_fifo))) = '1'), niosII_system_burst_4_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_4_upstream_waits_for_read) AND niosII_system_burst_4_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_4_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_4_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_4_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_4_upstream_transaction_burst_count, niosII_system_burst_4_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_4_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_4_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_4_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_4_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_4_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_4_upstream_current_burst <= niosII_system_burst_4_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_4_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_4_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_4_upstream_waits_for_read)) AND niosII_system_burst_4_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_4_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_4_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_4_upstream_waits_for_read)) AND NOT niosII_system_burst_4_upstream_load_fifo) OR niosII_system_burst_4_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_4_upstream_load_fifo <= p0_niosII_system_burst_4_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_4_upstream, which is an e_assign
  niosII_system_burst_4_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_4_upstream_current_burst_minus_one)) AND niosII_system_burst_4_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_4_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_4_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_4_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_4_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_4_upstream,
      full => open,
      clear_fifo => module_input99,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_4_upstream,
      read => niosII_system_burst_4_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input100,
      write => module_input101
    );

  module_input99 <= std_logic'('0');
  module_input100 <= std_logic'('0');
  module_input101 <= in_a_read_cycle AND NOT niosII_system_burst_4_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_4_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_4_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_4_upstream <= niosII_system_burst_4_upstream_readdatavalid_from_sa;
  --niosII_system_burst_4_upstream_writedata mux, which is an e_mux
  niosII_system_burst_4_upstream_writedata <= cpu_data_master_writedata;
  --byteaddress mux for niosII_system_burst_4/upstream, which is an e_mux
  niosII_system_burst_4_upstream_byteaddress <= cpu_data_master_address_to_slave (4 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_4_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_4_upstream;
  --cpu/data_master saved-grant niosII_system_burst_4/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_4_upstream <= internal_cpu_data_master_requests_niosII_system_burst_4_upstream;
  --allow new arb cycle for niosII_system_burst_4/upstream, which is an e_assign
  niosII_system_burst_4_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_4_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_4_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_4_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_4_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_4_upstream_begins_xfer) = '1'), niosII_system_burst_4_upstream_unreg_firsttransfer, niosII_system_burst_4_upstream_reg_firsttransfer);
  --niosII_system_burst_4_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_4_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_4_upstream_slavearbiterlockenable AND niosII_system_burst_4_upstream_any_continuerequest));
  --niosII_system_burst_4_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_4_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_4_upstream_begins_xfer) = '1' then 
        niosII_system_burst_4_upstream_reg_firsttransfer <= niosII_system_burst_4_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_4_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_4_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_4_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_4_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_4_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_4_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_4_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_4_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_4_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_4_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_4_upstream_begins_xfer) = '1' then 
        niosII_system_burst_4_upstream_bbt_burstcounter <= niosII_system_burst_4_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_4_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_4_upstream_beginbursttransfer_internal <= niosII_system_burst_4_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_4_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_4_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_4_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_4_upstream AND cpu_data_master_read;
  --niosII_system_burst_4_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_4_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_4_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_4_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_4_upstream_address mux, which is an e_mux
  niosII_system_burst_4_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_4_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_niosII_system_burst_4_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_4_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_4_upstream_end_xfer <= niosII_system_burst_4_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_4_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_4_upstream_waits_for_read <= niosII_system_burst_4_upstream_in_a_read_cycle AND internal_niosII_system_burst_4_upstream_waitrequest_from_sa;
  --niosII_system_burst_4_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_4_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_4_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_4_upstream_in_a_read_cycle;
  --niosII_system_burst_4_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_4_upstream_waits_for_write <= niosII_system_burst_4_upstream_in_a_write_cycle AND internal_niosII_system_burst_4_upstream_waitrequest_from_sa;
  --niosII_system_burst_4_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_4_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_4_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_4_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_4_upstream_counter <= std_logic'('0');
  --niosII_system_burst_4_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_4_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_4_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_4_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_4_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_4_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_4_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_4_upstream <= internal_cpu_data_master_granted_niosII_system_burst_4_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_4_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_4_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_4_upstream <= internal_cpu_data_master_requests_niosII_system_burst_4_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_4_upstream_burstcount <= internal_niosII_system_burst_4_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_4_upstream_read <= internal_niosII_system_burst_4_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_4_upstream_waitrequest_from_sa <= internal_niosII_system_burst_4_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_4_upstream_write <= internal_niosII_system_burst_4_upstream_write;
--synthesis translate_off
    --niosII_system_burst_4/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line143 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_4_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line143, now);
          write(write_line143, string'(": "));
          write(write_line143, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_4/upstream"));
          write(output, write_line143.all);
          deallocate (write_line143);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_4_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_4_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_4_downstream_granted_sysid_control_slave : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_qualified_request_sysid_control_slave : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_requests_sysid_control_slave : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal niosII_system_burst_4_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_4_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_4_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_4_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_4_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_4_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_4_downstream_arbitrator;


architecture europa of niosII_system_burst_4_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_4_downstream_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_niosII_system_burst_4_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_address_last_time :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_4_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_4_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_flush_niosII_system_burst_4_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_4_downstream_qualified_request_sysid_control_slave OR NOT niosII_system_burst_4_downstream_requests_sysid_control_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_4_downstream_qualified_request_sysid_control_slave OR NOT niosII_system_burst_4_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sysid_control_slave_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_4_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_4_downstream_qualified_request_sysid_control_slave OR NOT niosII_system_burst_4_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_4_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_4_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_4_downstream_address_to_slave <= niosII_system_burst_4_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_4_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_4_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_4_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave)))));
  --niosII_system_burst_4/downstream readdata mux, which is an e_mux
  niosII_system_burst_4_downstream_readdata <= sysid_control_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_4_downstream_waitrequest <= NOT niosII_system_burst_4_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_4_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_4_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_4_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_4_downstream_address_to_slave <= internal_niosII_system_burst_4_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_4_downstream_waitrequest <= internal_niosII_system_burst_4_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_4_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_4_downstream_address_last_time <= std_logic_vector'("000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_4_downstream_address_last_time <= niosII_system_burst_4_downstream_address;
      end if;

    end process;

    --niosII_system_burst_4/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_4_downstream_waitrequest AND ((niosII_system_burst_4_downstream_read OR niosII_system_burst_4_downstream_write));
      end if;

    end process;

    --niosII_system_burst_4_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line144 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_4_downstream_address /= niosII_system_burst_4_downstream_address_last_time))))) = '1' then 
          write(write_line144, now);
          write(write_line144, string'(": "));
          write(write_line144, string'("niosII_system_burst_4_downstream_address did not heed wait!!!"));
          write(output, write_line144.all);
          deallocate (write_line144);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_4_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_4_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_4_downstream_burstcount_last_time <= niosII_system_burst_4_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_4_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line145 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_4_downstream_burstcount) /= std_logic'(niosII_system_burst_4_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line145, now);
          write(write_line145, string'(": "));
          write(write_line145, string'("niosII_system_burst_4_downstream_burstcount did not heed wait!!!"));
          write(output, write_line145.all);
          deallocate (write_line145);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_4_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_4_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_4_downstream_byteenable_last_time <= niosII_system_burst_4_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_4_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line146 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_4_downstream_byteenable /= niosII_system_burst_4_downstream_byteenable_last_time))))) = '1' then 
          write(write_line146, now);
          write(write_line146, string'(": "));
          write(write_line146, string'("niosII_system_burst_4_downstream_byteenable did not heed wait!!!"));
          write(output, write_line146.all);
          deallocate (write_line146);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_4_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_4_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_4_downstream_read_last_time <= niosII_system_burst_4_downstream_read;
      end if;

    end process;

    --niosII_system_burst_4_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line147 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_4_downstream_read) /= std_logic'(niosII_system_burst_4_downstream_read_last_time)))))) = '1' then 
          write(write_line147, now);
          write(write_line147, string'(": "));
          write(write_line147, string'("niosII_system_burst_4_downstream_read did not heed wait!!!"));
          write(output, write_line147.all);
          deallocate (write_line147);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_4_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_4_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_4_downstream_write_last_time <= niosII_system_burst_4_downstream_write;
      end if;

    end process;

    --niosII_system_burst_4_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line148 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_4_downstream_write) /= std_logic'(niosII_system_burst_4_downstream_write_last_time)))))) = '1' then 
          write(write_line148, now);
          write(write_line148, string'(": "));
          write(write_line148, string'("niosII_system_burst_4_downstream_write did not heed wait!!!"));
          write(output, write_line148.all);
          deallocate (write_line148);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_4_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_4_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_4_downstream_writedata_last_time <= niosII_system_burst_4_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_4_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line149 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_4_downstream_writedata /= niosII_system_burst_4_downstream_writedata_last_time)))) AND niosII_system_burst_4_downstream_write)) = '1' then 
          write(write_line149, now);
          write(write_line149, string'(": "));
          write(write_line149, string'("niosII_system_burst_4_downstream_writedata did not heed wait!!!"));
          write(output, write_line149.all);
          deallocate (write_line149);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_5_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_5_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_5_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_5_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_5_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_5_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_5_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_5_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_5_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_5_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_5_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_5_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_5_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_5_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_5_upstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_5_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_5_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_5_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_5_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_5_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_5_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_5_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_5_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_5_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity niosII_system_burst_5_upstream_arbitrator;


architecture europa of niosII_system_burst_5_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_5_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_5_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_5_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_5_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_5_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_5_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_5_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_5_upstream_write :  STD_LOGIC;
                signal module_input102 :  STD_LOGIC;
                signal module_input103 :  STD_LOGIC;
                signal module_input104 :  STD_LOGIC;
                signal module_input105 :  STD_LOGIC;
                signal module_input106 :  STD_LOGIC;
                signal module_input107 :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_5_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_5_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_5_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_5_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_5_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_5_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_5_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_5_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_5_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_5_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_5_upstream);
  --assign niosII_system_burst_5_upstream_readdatavalid_from_sa = niosII_system_burst_5_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_5_upstream_readdatavalid_from_sa <= niosII_system_burst_5_upstream_readdatavalid;
  --assign niosII_system_burst_5_upstream_readdata_from_sa = niosII_system_burst_5_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_5_upstream_readdata_from_sa <= niosII_system_burst_5_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_5_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1100100001001000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_5_upstream_waitrequest_from_sa = niosII_system_burst_5_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_5_upstream_waitrequest_from_sa <= niosII_system_burst_5_upstream_waitrequest;
  --niosII_system_burst_5_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_5_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_5_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_5_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_5_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_5_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_5_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_5_upstream;
  --niosII_system_burst_5_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_5_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_5_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_5_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_5_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_5_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_5_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_5_upstream_allgrants <= niosII_system_burst_5_upstream_grant_vector;
  --niosII_system_burst_5_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_5_upstream_end_xfer <= NOT ((niosII_system_burst_5_upstream_waits_for_read OR niosII_system_burst_5_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_5_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_5_upstream <= niosII_system_burst_5_upstream_end_xfer AND (((NOT niosII_system_burst_5_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_5_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_5_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_5_upstream AND niosII_system_burst_5_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_5_upstream AND NOT niosII_system_burst_5_upstream_non_bursting_master_requests));
  --niosII_system_burst_5_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_5_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_5_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_5_upstream_arb_share_counter <= niosII_system_burst_5_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_5_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_5_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_5_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_5_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_5_upstream AND NOT niosII_system_burst_5_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_5_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_5_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_5/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_5_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_5_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_5_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_5_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_5/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_5_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_5_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_5_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_5_upstream <= internal_cpu_data_master_requests_niosII_system_burst_5_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_5_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_5_upstream_move_on_to_next_transaction <= niosII_system_burst_5_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_5_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_5_upstream, which is an e_mux
  niosII_system_burst_5_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_5_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_5_upstream : burstcount_fifo_for_niosII_system_burst_5_upstream_module
    port map(
      data_out => niosII_system_burst_5_upstream_transaction_burst_count,
      empty => niosII_system_burst_5_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input102,
      clk => clk,
      data_in => niosII_system_burst_5_upstream_selected_burstcount,
      read => niosII_system_burst_5_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input103,
      write => module_input104
    );

  module_input102 <= std_logic'('0');
  module_input103 <= std_logic'('0');
  module_input104 <= ((in_a_read_cycle AND NOT niosII_system_burst_5_upstream_waits_for_read) AND niosII_system_burst_5_upstream_load_fifo) AND NOT ((niosII_system_burst_5_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_5_upstream_burstcount_fifo_empty));

  --niosII_system_burst_5_upstream current burst minus one, which is an e_assign
  niosII_system_burst_5_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_5_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_5_upstream, which is an e_mux
  niosII_system_burst_5_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_5_upstream_waits_for_read)) AND NOT niosII_system_burst_5_upstream_load_fifo))) = '1'), niosII_system_burst_5_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_5_upstream_waits_for_read) AND niosII_system_burst_5_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_5_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_5_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_5_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_5_upstream_transaction_burst_count, niosII_system_burst_5_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_5_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_5_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_5_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_5_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_5_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_5_upstream_current_burst <= niosII_system_burst_5_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_5_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_5_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_5_upstream_waits_for_read)) AND niosII_system_burst_5_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_5_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_5_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_5_upstream_waits_for_read)) AND NOT niosII_system_burst_5_upstream_load_fifo) OR niosII_system_burst_5_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_5_upstream_load_fifo <= p0_niosII_system_burst_5_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_5_upstream, which is an e_assign
  niosII_system_burst_5_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_5_upstream_current_burst_minus_one)) AND niosII_system_burst_5_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_5_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_5_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_5_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_5_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_5_upstream,
      full => open,
      clear_fifo => module_input105,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_5_upstream,
      read => niosII_system_burst_5_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input106,
      write => module_input107
    );

  module_input105 <= std_logic'('0');
  module_input106 <= std_logic'('0');
  module_input107 <= in_a_read_cycle AND NOT niosII_system_burst_5_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_5_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_5_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_5_upstream <= niosII_system_burst_5_upstream_readdatavalid_from_sa;
  --niosII_system_burst_5_upstream_writedata mux, which is an e_mux
  niosII_system_burst_5_upstream_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --byteaddress mux for niosII_system_burst_5/upstream, which is an e_mux
  niosII_system_burst_5_upstream_byteaddress <= cpu_data_master_address_to_slave (4 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_5_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_5_upstream;
  --cpu/data_master saved-grant niosII_system_burst_5/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_5_upstream <= internal_cpu_data_master_requests_niosII_system_burst_5_upstream;
  --allow new arb cycle for niosII_system_burst_5/upstream, which is an e_assign
  niosII_system_burst_5_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_5_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_5_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_5_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_5_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_5_upstream_begins_xfer) = '1'), niosII_system_burst_5_upstream_unreg_firsttransfer, niosII_system_burst_5_upstream_reg_firsttransfer);
  --niosII_system_burst_5_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_5_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_5_upstream_slavearbiterlockenable AND niosII_system_burst_5_upstream_any_continuerequest));
  --niosII_system_burst_5_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_5_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_5_upstream_begins_xfer) = '1' then 
        niosII_system_burst_5_upstream_reg_firsttransfer <= niosII_system_burst_5_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_5_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_5_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_5_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_5_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_5_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_5_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_5_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_5_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_5_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_5_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_5_upstream_begins_xfer) = '1' then 
        niosII_system_burst_5_upstream_bbt_burstcounter <= niosII_system_burst_5_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_5_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_5_upstream_beginbursttransfer_internal <= niosII_system_burst_5_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_5_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_5_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_5_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_5_upstream AND cpu_data_master_read;
  --niosII_system_burst_5_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_5_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_5_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_5_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_5_upstream_address mux, which is an e_mux
  niosII_system_burst_5_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_5_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --d1_niosII_system_burst_5_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_5_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_5_upstream_end_xfer <= niosII_system_burst_5_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_5_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_5_upstream_waits_for_read <= niosII_system_burst_5_upstream_in_a_read_cycle AND internal_niosII_system_burst_5_upstream_waitrequest_from_sa;
  --niosII_system_burst_5_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_5_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_5_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_5_upstream_in_a_read_cycle;
  --niosII_system_burst_5_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_5_upstream_waits_for_write <= niosII_system_burst_5_upstream_in_a_write_cycle AND internal_niosII_system_burst_5_upstream_waitrequest_from_sa;
  --niosII_system_burst_5_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_5_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_5_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_5_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_5_upstream_counter <= std_logic'('0');
  --niosII_system_burst_5_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_5_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_5_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_5_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_5_upstream <= internal_cpu_data_master_granted_niosII_system_burst_5_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_5_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_5_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_5_upstream <= internal_cpu_data_master_requests_niosII_system_burst_5_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_5_upstream_burstcount <= internal_niosII_system_burst_5_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_5_upstream_read <= internal_niosII_system_burst_5_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_5_upstream_waitrequest_from_sa <= internal_niosII_system_burst_5_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_5_upstream_write <= internal_niosII_system_burst_5_upstream_write;
--synthesis translate_off
    --niosII_system_burst_5/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line150 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_5_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line150, now);
          write(write_line150, string'(": "));
          write(write_line150, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_5/upstream"));
          write(output, write_line150.all);
          deallocate (write_line150);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_5_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sys_clk_timer_s1_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_5_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal niosII_system_burst_5_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_5_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_5_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_5_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_5_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_5_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_5_downstream_arbitrator;


architecture europa of niosII_system_burst_5_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_5_downstream_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_5_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_5_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_flush_niosII_system_burst_5_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 OR NOT niosII_system_burst_5_downstream_requests_sys_clk_timer_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 OR NOT niosII_system_burst_5_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sys_clk_timer_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_5_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 OR NOT niosII_system_burst_5_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_5_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_5_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_5_downstream_address_to_slave <= niosII_system_burst_5_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_5_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_5_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_5_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1)))));
  --niosII_system_burst_5/downstream readdata mux, which is an e_mux
  niosII_system_burst_5_downstream_readdata <= sys_clk_timer_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_5_downstream_waitrequest <= NOT niosII_system_burst_5_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_5_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_5_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_5_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_5_downstream_address_to_slave <= internal_niosII_system_burst_5_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_5_downstream_waitrequest <= internal_niosII_system_burst_5_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_5_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_5_downstream_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_5_downstream_address_last_time <= niosII_system_burst_5_downstream_address;
      end if;

    end process;

    --niosII_system_burst_5/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_5_downstream_waitrequest AND ((niosII_system_burst_5_downstream_read OR niosII_system_burst_5_downstream_write));
      end if;

    end process;

    --niosII_system_burst_5_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line151 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_5_downstream_address /= niosII_system_burst_5_downstream_address_last_time))))) = '1' then 
          write(write_line151, now);
          write(write_line151, string'(": "));
          write(write_line151, string'("niosII_system_burst_5_downstream_address did not heed wait!!!"));
          write(output, write_line151.all);
          deallocate (write_line151);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_5_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_5_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_5_downstream_burstcount_last_time <= niosII_system_burst_5_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_5_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line152 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_5_downstream_burstcount) /= std_logic'(niosII_system_burst_5_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line152, now);
          write(write_line152, string'(": "));
          write(write_line152, string'("niosII_system_burst_5_downstream_burstcount did not heed wait!!!"));
          write(output, write_line152.all);
          deallocate (write_line152);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_5_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_5_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_5_downstream_byteenable_last_time <= niosII_system_burst_5_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_5_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line153 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_5_downstream_byteenable /= niosII_system_burst_5_downstream_byteenable_last_time))))) = '1' then 
          write(write_line153, now);
          write(write_line153, string'(": "));
          write(write_line153, string'("niosII_system_burst_5_downstream_byteenable did not heed wait!!!"));
          write(output, write_line153.all);
          deallocate (write_line153);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_5_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_5_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_5_downstream_read_last_time <= niosII_system_burst_5_downstream_read;
      end if;

    end process;

    --niosII_system_burst_5_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line154 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_5_downstream_read) /= std_logic'(niosII_system_burst_5_downstream_read_last_time)))))) = '1' then 
          write(write_line154, now);
          write(write_line154, string'(": "));
          write(write_line154, string'("niosII_system_burst_5_downstream_read did not heed wait!!!"));
          write(output, write_line154.all);
          deallocate (write_line154);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_5_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_5_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_5_downstream_write_last_time <= niosII_system_burst_5_downstream_write;
      end if;

    end process;

    --niosII_system_burst_5_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line155 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_5_downstream_write) /= std_logic'(niosII_system_burst_5_downstream_write_last_time)))))) = '1' then 
          write(write_line155, now);
          write(write_line155, string'(": "));
          write(write_line155, string'("niosII_system_burst_5_downstream_write did not heed wait!!!"));
          write(output, write_line155.all);
          deallocate (write_line155);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_5_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_5_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_5_downstream_writedata_last_time <= niosII_system_burst_5_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_5_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line156 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_5_downstream_writedata /= niosII_system_burst_5_downstream_writedata_last_time)))) AND niosII_system_burst_5_downstream_write)) = '1' then 
          write(write_line156, now);
          write(write_line156, string'(": "));
          write(write_line156, string'("niosII_system_burst_5_downstream_writedata did not heed wait!!!"));
          write(output, write_line156.all);
          deallocate (write_line156);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_6_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_6_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_6_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_6_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_6_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_6_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_6_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_6_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_6_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_6_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_6_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_6_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_6_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_6_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_6_upstream_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_6_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_6_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_6_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_6_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_6_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_6_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_6_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_6_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_6_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity niosII_system_burst_6_upstream_arbitrator;


architecture europa of niosII_system_burst_6_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_6_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_6_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_6_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_6_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_6_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_6_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_6_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_6_upstream_write :  STD_LOGIC;
                signal module_input108 :  STD_LOGIC;
                signal module_input109 :  STD_LOGIC;
                signal module_input110 :  STD_LOGIC;
                signal module_input111 :  STD_LOGIC;
                signal module_input112 :  STD_LOGIC;
                signal module_input113 :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_6_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_6_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_6_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_6_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_6_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_6_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_6_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_6_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_6_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_6_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_6_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_6_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_6_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_6_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_6_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_6_upstream);
  --assign niosII_system_burst_6_upstream_readdatavalid_from_sa = niosII_system_burst_6_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_6_upstream_readdatavalid_from_sa <= niosII_system_burst_6_upstream_readdatavalid;
  --assign niosII_system_burst_6_upstream_readdata_from_sa = niosII_system_burst_6_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_6_upstream_readdata_from_sa <= niosII_system_burst_6_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_6_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("1100100001001000011011000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_6_upstream_waitrequest_from_sa = niosII_system_burst_6_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_6_upstream_waitrequest_from_sa <= niosII_system_burst_6_upstream_waitrequest;
  --niosII_system_burst_6_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_6_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_6_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_6_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_6_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_6_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_6_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_6_upstream;
  --niosII_system_burst_6_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_6_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_6_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_6_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_6_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_6_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_6_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_6_upstream_allgrants <= niosII_system_burst_6_upstream_grant_vector;
  --niosII_system_burst_6_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_6_upstream_end_xfer <= NOT ((niosII_system_burst_6_upstream_waits_for_read OR niosII_system_burst_6_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_6_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_6_upstream <= niosII_system_burst_6_upstream_end_xfer AND (((NOT niosII_system_burst_6_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_6_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_6_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_6_upstream AND niosII_system_burst_6_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_6_upstream AND NOT niosII_system_burst_6_upstream_non_bursting_master_requests));
  --niosII_system_burst_6_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_6_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_6_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_6_upstream_arb_share_counter <= niosII_system_burst_6_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_6_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_6_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_6_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_6_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_6_upstream AND NOT niosII_system_burst_6_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_6_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_6_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_6/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_6_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_6_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_6_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_6_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_6/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_6_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_6_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_6_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_6_upstream <= internal_cpu_data_master_requests_niosII_system_burst_6_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_6_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_6_upstream_move_on_to_next_transaction <= niosII_system_burst_6_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_6_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_6_upstream, which is an e_mux
  niosII_system_burst_6_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_6_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_6_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_6_upstream : burstcount_fifo_for_niosII_system_burst_6_upstream_module
    port map(
      data_out => niosII_system_burst_6_upstream_transaction_burst_count,
      empty => niosII_system_burst_6_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input108,
      clk => clk,
      data_in => niosII_system_burst_6_upstream_selected_burstcount,
      read => niosII_system_burst_6_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input109,
      write => module_input110
    );

  module_input108 <= std_logic'('0');
  module_input109 <= std_logic'('0');
  module_input110 <= ((in_a_read_cycle AND NOT niosII_system_burst_6_upstream_waits_for_read) AND niosII_system_burst_6_upstream_load_fifo) AND NOT ((niosII_system_burst_6_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_6_upstream_burstcount_fifo_empty));

  --niosII_system_burst_6_upstream current burst minus one, which is an e_assign
  niosII_system_burst_6_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_6_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_6_upstream, which is an e_mux
  niosII_system_burst_6_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_6_upstream_waits_for_read)) AND NOT niosII_system_burst_6_upstream_load_fifo))) = '1'), niosII_system_burst_6_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_6_upstream_waits_for_read) AND niosII_system_burst_6_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_6_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_6_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_6_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_6_upstream_transaction_burst_count, niosII_system_burst_6_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_6_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_6_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_6_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_6_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_6_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_6_upstream_current_burst <= niosII_system_burst_6_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_6_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_6_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_6_upstream_waits_for_read)) AND niosII_system_burst_6_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_6_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_6_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_6_upstream_waits_for_read)) AND NOT niosII_system_burst_6_upstream_load_fifo) OR niosII_system_burst_6_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_6_upstream_load_fifo <= p0_niosII_system_burst_6_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_6_upstream, which is an e_assign
  niosII_system_burst_6_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_6_upstream_current_burst_minus_one)) AND niosII_system_burst_6_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_6_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_6_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_6_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_6_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_6_upstream,
      full => open,
      clear_fifo => module_input111,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_6_upstream,
      read => niosII_system_burst_6_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input112,
      write => module_input113
    );

  module_input111 <= std_logic'('0');
  module_input112 <= std_logic'('0');
  module_input113 <= in_a_read_cycle AND NOT niosII_system_burst_6_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_6_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_6_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_6_upstream <= niosII_system_burst_6_upstream_readdatavalid_from_sa;
  --niosII_system_burst_6_upstream_writedata mux, which is an e_mux
  niosII_system_burst_6_upstream_writedata <= cpu_data_master_writedata;
  --byteaddress mux for niosII_system_burst_6/upstream, which is an e_mux
  niosII_system_burst_6_upstream_byteaddress <= cpu_data_master_address_to_slave (4 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_6_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_6_upstream;
  --cpu/data_master saved-grant niosII_system_burst_6/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_6_upstream <= internal_cpu_data_master_requests_niosII_system_burst_6_upstream;
  --allow new arb cycle for niosII_system_burst_6/upstream, which is an e_assign
  niosII_system_burst_6_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_6_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_6_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_6_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_6_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_6_upstream_begins_xfer) = '1'), niosII_system_burst_6_upstream_unreg_firsttransfer, niosII_system_burst_6_upstream_reg_firsttransfer);
  --niosII_system_burst_6_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_6_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_6_upstream_slavearbiterlockenable AND niosII_system_burst_6_upstream_any_continuerequest));
  --niosII_system_burst_6_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_6_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_6_upstream_begins_xfer) = '1' then 
        niosII_system_burst_6_upstream_reg_firsttransfer <= niosII_system_burst_6_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_6_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_6_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_6_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_6_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_6_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_6_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_6_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_6_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_6_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_6_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_6_upstream_begins_xfer) = '1' then 
        niosII_system_burst_6_upstream_bbt_burstcounter <= niosII_system_burst_6_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_6_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_6_upstream_beginbursttransfer_internal <= niosII_system_burst_6_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_6_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_6_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_6_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_6_upstream AND cpu_data_master_read;
  --niosII_system_burst_6_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_6_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_6_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_6_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_6_upstream_address mux, which is an e_mux
  niosII_system_burst_6_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_6_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_niosII_system_burst_6_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_6_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_6_upstream_end_xfer <= niosII_system_burst_6_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_6_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_6_upstream_waits_for_read <= niosII_system_burst_6_upstream_in_a_read_cycle AND internal_niosII_system_burst_6_upstream_waitrequest_from_sa;
  --niosII_system_burst_6_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_6_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_6_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_6_upstream_in_a_read_cycle;
  --niosII_system_burst_6_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_6_upstream_waits_for_write <= niosII_system_burst_6_upstream_in_a_write_cycle AND internal_niosII_system_burst_6_upstream_waitrequest_from_sa;
  --niosII_system_burst_6_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_6_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_6_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_6_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_6_upstream_counter <= std_logic'('0');
  --niosII_system_burst_6_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_6_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_6_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_6_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_6_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_6_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_6_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_6_upstream <= internal_cpu_data_master_granted_niosII_system_burst_6_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_6_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_6_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_6_upstream <= internal_cpu_data_master_requests_niosII_system_burst_6_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_6_upstream_burstcount <= internal_niosII_system_burst_6_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_6_upstream_read <= internal_niosII_system_burst_6_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_6_upstream_waitrequest_from_sa <= internal_niosII_system_burst_6_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_6_upstream_write <= internal_niosII_system_burst_6_upstream_write;
--synthesis translate_off
    --niosII_system_burst_6/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line157 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_6_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line157, now);
          write(write_line157, string'(": "));
          write(write_line157, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_6/upstream"));
          write(output, write_line157.all);
          deallocate (write_line157);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_6_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_6_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_6_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_6_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_6_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_6_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_6_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_6_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_6_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_6_downstream_arbitrator;


architecture europa of niosII_system_burst_6_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_6_downstream_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_niosII_system_burst_6_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_address_last_time :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_6_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_6_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_flush_niosII_system_burst_6_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave OR NOT niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave OR NOT ((niosII_system_burst_6_downstream_read OR niosII_system_burst_6_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_6_downstream_read OR niosII_system_burst_6_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave OR NOT ((niosII_system_burst_6_downstream_read OR niosII_system_burst_6_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_6_downstream_read OR niosII_system_burst_6_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_6_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_6_downstream_address_to_slave <= niosII_system_burst_6_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_6_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_6_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_6_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave)))));
  --niosII_system_burst_6/downstream readdata mux, which is an e_mux
  niosII_system_burst_6_downstream_readdata <= jtag_uart_avalon_jtag_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_6_downstream_waitrequest <= NOT niosII_system_burst_6_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_6_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_6_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_6_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_6_downstream_address_to_slave <= internal_niosII_system_burst_6_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_6_downstream_waitrequest <= internal_niosII_system_burst_6_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_6_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_6_downstream_address_last_time <= std_logic_vector'("000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_6_downstream_address_last_time <= niosII_system_burst_6_downstream_address;
      end if;

    end process;

    --niosII_system_burst_6/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_6_downstream_waitrequest AND ((niosII_system_burst_6_downstream_read OR niosII_system_burst_6_downstream_write));
      end if;

    end process;

    --niosII_system_burst_6_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line158 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_6_downstream_address /= niosII_system_burst_6_downstream_address_last_time))))) = '1' then 
          write(write_line158, now);
          write(write_line158, string'(": "));
          write(write_line158, string'("niosII_system_burst_6_downstream_address did not heed wait!!!"));
          write(output, write_line158.all);
          deallocate (write_line158);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_6_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_6_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_6_downstream_burstcount_last_time <= niosII_system_burst_6_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_6_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line159 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_6_downstream_burstcount) /= std_logic'(niosII_system_burst_6_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line159, now);
          write(write_line159, string'(": "));
          write(write_line159, string'("niosII_system_burst_6_downstream_burstcount did not heed wait!!!"));
          write(output, write_line159.all);
          deallocate (write_line159);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_6_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_6_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_6_downstream_byteenable_last_time <= niosII_system_burst_6_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_6_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line160 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_6_downstream_byteenable /= niosII_system_burst_6_downstream_byteenable_last_time))))) = '1' then 
          write(write_line160, now);
          write(write_line160, string'(": "));
          write(write_line160, string'("niosII_system_burst_6_downstream_byteenable did not heed wait!!!"));
          write(output, write_line160.all);
          deallocate (write_line160);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_6_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_6_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_6_downstream_read_last_time <= niosII_system_burst_6_downstream_read;
      end if;

    end process;

    --niosII_system_burst_6_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line161 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_6_downstream_read) /= std_logic'(niosII_system_burst_6_downstream_read_last_time)))))) = '1' then 
          write(write_line161, now);
          write(write_line161, string'(": "));
          write(write_line161, string'("niosII_system_burst_6_downstream_read did not heed wait!!!"));
          write(output, write_line161.all);
          deallocate (write_line161);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_6_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_6_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_6_downstream_write_last_time <= niosII_system_burst_6_downstream_write;
      end if;

    end process;

    --niosII_system_burst_6_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line162 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_6_downstream_write) /= std_logic'(niosII_system_burst_6_downstream_write_last_time)))))) = '1' then 
          write(write_line162, now);
          write(write_line162, string'(": "));
          write(write_line162, string'("niosII_system_burst_6_downstream_write did not heed wait!!!"));
          write(output, write_line162.all);
          deallocate (write_line162);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_6_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_6_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_6_downstream_writedata_last_time <= niosII_system_burst_6_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_6_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line163 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_6_downstream_writedata /= niosII_system_burst_6_downstream_writedata_last_time)))) AND niosII_system_burst_6_downstream_write)) = '1' then 
          write(write_line163, now);
          write(write_line163, string'(": "));
          write(write_line163, string'("niosII_system_burst_6_downstream_writedata did not heed wait!!!"));
          write(output, write_line163.all);
          deallocate (write_line163);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_7_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_7_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_7_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_7_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_7_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_7_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_7_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_7_upstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_7_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_7_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_7_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_7_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_7_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_7_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_7_upstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_7_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_7_upstream_byteaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_7_upstream_byteenable : OUT STD_LOGIC;
                 signal niosII_system_burst_7_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_7_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_7_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_7_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_7_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_7_upstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity niosII_system_burst_7_upstream_arbitrator;


architecture europa of niosII_system_burst_7_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_7_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_7_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_7_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_7_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_7_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_7_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_7_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_7_upstream_write :  STD_LOGIC;
                signal module_input114 :  STD_LOGIC;
                signal module_input115 :  STD_LOGIC;
                signal module_input116 :  STD_LOGIC;
                signal module_input117 :  STD_LOGIC;
                signal module_input118 :  STD_LOGIC;
                signal module_input119 :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_7_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_7_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_7_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_7_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_7_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_7_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_7_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_7_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_7_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_7_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_7_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_7_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_7_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_7_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_7_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_7_upstream);
  --assign niosII_system_burst_7_upstream_readdatavalid_from_sa = niosII_system_burst_7_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_7_upstream_readdatavalid_from_sa <= niosII_system_burst_7_upstream_readdatavalid;
  --assign niosII_system_burst_7_upstream_readdata_from_sa = niosII_system_burst_7_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_7_upstream_readdata_from_sa <= niosII_system_burst_7_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_7_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1100100001001000010000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_7_upstream_waitrequest_from_sa = niosII_system_burst_7_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_7_upstream_waitrequest_from_sa <= niosII_system_burst_7_upstream_waitrequest;
  --niosII_system_burst_7_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_7_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_7_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_7_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_7_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_7_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_7_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_7_upstream;
  --niosII_system_burst_7_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_7_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_7_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_7_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_7_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_7_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_7_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_7_upstream_allgrants <= niosII_system_burst_7_upstream_grant_vector;
  --niosII_system_burst_7_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_7_upstream_end_xfer <= NOT ((niosII_system_burst_7_upstream_waits_for_read OR niosII_system_burst_7_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_7_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_7_upstream <= niosII_system_burst_7_upstream_end_xfer AND (((NOT niosII_system_burst_7_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_7_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_7_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_7_upstream AND niosII_system_burst_7_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_7_upstream AND NOT niosII_system_burst_7_upstream_non_bursting_master_requests));
  --niosII_system_burst_7_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_7_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_7_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_7_upstream_arb_share_counter <= niosII_system_burst_7_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_7_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_7_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_7_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_7_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_7_upstream AND NOT niosII_system_burst_7_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_7_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_7_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_7/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_7_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_7_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_7_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_7_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_7/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_7_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_7_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_7_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_7_upstream <= internal_cpu_data_master_requests_niosII_system_burst_7_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_7_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_7_upstream_move_on_to_next_transaction <= niosII_system_burst_7_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_7_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_7_upstream, which is an e_mux
  niosII_system_burst_7_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_7_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_7_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_7_upstream : burstcount_fifo_for_niosII_system_burst_7_upstream_module
    port map(
      data_out => niosII_system_burst_7_upstream_transaction_burst_count,
      empty => niosII_system_burst_7_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input114,
      clk => clk,
      data_in => niosII_system_burst_7_upstream_selected_burstcount,
      read => niosII_system_burst_7_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input115,
      write => module_input116
    );

  module_input114 <= std_logic'('0');
  module_input115 <= std_logic'('0');
  module_input116 <= ((in_a_read_cycle AND NOT niosII_system_burst_7_upstream_waits_for_read) AND niosII_system_burst_7_upstream_load_fifo) AND NOT ((niosII_system_burst_7_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_7_upstream_burstcount_fifo_empty));

  --niosII_system_burst_7_upstream current burst minus one, which is an e_assign
  niosII_system_burst_7_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_7_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_7_upstream, which is an e_mux
  niosII_system_burst_7_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_7_upstream_waits_for_read)) AND NOT niosII_system_burst_7_upstream_load_fifo))) = '1'), niosII_system_burst_7_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_7_upstream_waits_for_read) AND niosII_system_burst_7_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_7_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_7_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_7_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_7_upstream_transaction_burst_count, niosII_system_burst_7_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_7_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_7_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_7_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_7_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_7_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_7_upstream_current_burst <= niosII_system_burst_7_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_7_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_7_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_7_upstream_waits_for_read)) AND niosII_system_burst_7_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_7_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_7_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_7_upstream_waits_for_read)) AND NOT niosII_system_burst_7_upstream_load_fifo) OR niosII_system_burst_7_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_7_upstream_load_fifo <= p0_niosII_system_burst_7_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_7_upstream, which is an e_assign
  niosII_system_burst_7_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_7_upstream_current_burst_minus_one)) AND niosII_system_burst_7_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_7_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_7_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_7_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_7_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_7_upstream,
      full => open,
      clear_fifo => module_input117,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_7_upstream,
      read => niosII_system_burst_7_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input118,
      write => module_input119
    );

  module_input117 <= std_logic'('0');
  module_input118 <= std_logic'('0');
  module_input119 <= in_a_read_cycle AND NOT niosII_system_burst_7_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_7_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_7_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_7_upstream <= niosII_system_burst_7_upstream_readdatavalid_from_sa;
  --niosII_system_burst_7_upstream_writedata mux, which is an e_mux
  niosII_system_burst_7_upstream_writedata <= cpu_data_master_writedata (7 DOWNTO 0);
  --byteaddress mux for niosII_system_burst_7/upstream, which is an e_mux
  niosII_system_burst_7_upstream_byteaddress <= cpu_data_master_address_to_slave (1 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_7_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_7_upstream;
  --cpu/data_master saved-grant niosII_system_burst_7/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_7_upstream <= internal_cpu_data_master_requests_niosII_system_burst_7_upstream;
  --allow new arb cycle for niosII_system_burst_7/upstream, which is an e_assign
  niosII_system_burst_7_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_7_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_7_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_7_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_7_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_7_upstream_begins_xfer) = '1'), niosII_system_burst_7_upstream_unreg_firsttransfer, niosII_system_burst_7_upstream_reg_firsttransfer);
  --niosII_system_burst_7_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_7_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_7_upstream_slavearbiterlockenable AND niosII_system_burst_7_upstream_any_continuerequest));
  --niosII_system_burst_7_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_7_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_7_upstream_begins_xfer) = '1' then 
        niosII_system_burst_7_upstream_reg_firsttransfer <= niosII_system_burst_7_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_7_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_7_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_7_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_7_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_7_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_7_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_7_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_7_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_7_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_7_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_7_upstream_begins_xfer) = '1' then 
        niosII_system_burst_7_upstream_bbt_burstcounter <= niosII_system_burst_7_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_7_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_7_upstream_beginbursttransfer_internal <= niosII_system_burst_7_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_7_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_7_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_7_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_7_upstream AND cpu_data_master_read;
  --niosII_system_burst_7_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_7_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_7_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_7_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_7_upstream_address mux, which is an e_mux
  niosII_system_burst_7_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_7_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_niosII_system_burst_7_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_7_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_7_upstream_end_xfer <= niosII_system_burst_7_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_7_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_7_upstream_waits_for_read <= niosII_system_burst_7_upstream_in_a_read_cycle AND internal_niosII_system_burst_7_upstream_waitrequest_from_sa;
  --niosII_system_burst_7_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_7_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_7_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_7_upstream_in_a_read_cycle;
  --niosII_system_burst_7_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_7_upstream_waits_for_write <= niosII_system_burst_7_upstream_in_a_write_cycle AND internal_niosII_system_burst_7_upstream_waitrequest_from_sa;
  --niosII_system_burst_7_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_7_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_7_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_7_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_7_upstream_counter <= std_logic'('0');
  --niosII_system_burst_7_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_7_upstream_byteenable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_7_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_7_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_7_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_7_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_7_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_7_upstream <= internal_cpu_data_master_granted_niosII_system_burst_7_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_7_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_7_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_7_upstream <= internal_cpu_data_master_requests_niosII_system_burst_7_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_7_upstream_burstcount <= internal_niosII_system_burst_7_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_7_upstream_read <= internal_niosII_system_burst_7_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_7_upstream_waitrequest_from_sa <= internal_niosII_system_burst_7_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_7_upstream_write <= internal_niosII_system_burst_7_upstream_write;
--synthesis translate_off
    --niosII_system_burst_7/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line164 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_7_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line164, now);
          write(write_line164, string'(": "));
          write(write_line164, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_7/upstream"));
          write(output, write_line164.all);
          deallocate (write_line164);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_7_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_lcd_display_control_slave_end_xfer : IN STD_LOGIC;
                 signal lcd_display_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal lcd_display_control_slave_wait_counter_eq_0 : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_7_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_byteenable : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_granted_lcd_display_control_slave : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_requests_lcd_display_control_slave : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_7_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_7_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_7_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_7_downstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_7_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_7_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_7_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_7_downstream_arbitrator;


architecture europa of niosII_system_burst_7_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_7_downstream_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_niosII_system_burst_7_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_7_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_byteenable_last_time :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pre_flush_niosII_system_burst_7_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave OR NOT niosII_system_burst_7_downstream_requests_lcd_display_control_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave OR NOT niosII_system_burst_7_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((lcd_display_control_slave_wait_counter_eq_0 AND NOT d1_lcd_display_control_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_7_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave OR NOT niosII_system_burst_7_downstream_write)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((lcd_display_control_slave_wait_counter_eq_0 AND NOT d1_lcd_display_control_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_7_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_7_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_7_downstream_address_to_slave <= niosII_system_burst_7_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_7_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_7_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_7_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave)))));
  --niosII_system_burst_7/downstream readdata mux, which is an e_mux
  niosII_system_burst_7_downstream_readdata <= lcd_display_control_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_7_downstream_waitrequest <= NOT niosII_system_burst_7_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_7_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_7_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_7_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_7_downstream_address_to_slave <= internal_niosII_system_burst_7_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_7_downstream_waitrequest <= internal_niosII_system_burst_7_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_7_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_7_downstream_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_7_downstream_address_last_time <= niosII_system_burst_7_downstream_address;
      end if;

    end process;

    --niosII_system_burst_7/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_7_downstream_waitrequest AND ((niosII_system_burst_7_downstream_read OR niosII_system_burst_7_downstream_write));
      end if;

    end process;

    --niosII_system_burst_7_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line165 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_7_downstream_address /= niosII_system_burst_7_downstream_address_last_time))))) = '1' then 
          write(write_line165, now);
          write(write_line165, string'(": "));
          write(write_line165, string'("niosII_system_burst_7_downstream_address did not heed wait!!!"));
          write(output, write_line165.all);
          deallocate (write_line165);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_7_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_7_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_7_downstream_burstcount_last_time <= niosII_system_burst_7_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_7_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line166 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_7_downstream_burstcount) /= std_logic'(niosII_system_burst_7_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line166, now);
          write(write_line166, string'(": "));
          write(write_line166, string'("niosII_system_burst_7_downstream_burstcount did not heed wait!!!"));
          write(output, write_line166.all);
          deallocate (write_line166);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_7_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_7_downstream_byteenable_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_7_downstream_byteenable_last_time <= niosII_system_burst_7_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_7_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line167 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_7_downstream_byteenable) /= std_logic'(niosII_system_burst_7_downstream_byteenable_last_time)))))) = '1' then 
          write(write_line167, now);
          write(write_line167, string'(": "));
          write(write_line167, string'("niosII_system_burst_7_downstream_byteenable did not heed wait!!!"));
          write(output, write_line167.all);
          deallocate (write_line167);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_7_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_7_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_7_downstream_read_last_time <= niosII_system_burst_7_downstream_read;
      end if;

    end process;

    --niosII_system_burst_7_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line168 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_7_downstream_read) /= std_logic'(niosII_system_burst_7_downstream_read_last_time)))))) = '1' then 
          write(write_line168, now);
          write(write_line168, string'(": "));
          write(write_line168, string'("niosII_system_burst_7_downstream_read did not heed wait!!!"));
          write(output, write_line168.all);
          deallocate (write_line168);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_7_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_7_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_7_downstream_write_last_time <= niosII_system_burst_7_downstream_write;
      end if;

    end process;

    --niosII_system_burst_7_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line169 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_7_downstream_write) /= std_logic'(niosII_system_burst_7_downstream_write_last_time)))))) = '1' then 
          write(write_line169, now);
          write(write_line169, string'(": "));
          write(write_line169, string'("niosII_system_burst_7_downstream_write did not heed wait!!!"));
          write(output, write_line169.all);
          deallocate (write_line169);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_7_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_7_downstream_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_7_downstream_writedata_last_time <= niosII_system_burst_7_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_7_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line170 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_7_downstream_writedata /= niosII_system_burst_7_downstream_writedata_last_time)))) AND niosII_system_burst_7_downstream_write)) = '1' then 
          write(write_line170, now);
          write(write_line170, string'(": "));
          write(write_line170, string'("niosII_system_burst_7_downstream_writedata did not heed wait!!!"));
          write(output, write_line170.all);
          deallocate (write_line170);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_8_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_8_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_8_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_8_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_8_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_8_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_8_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_8_upstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_8_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_8_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_8_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_8_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_8_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_8_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_8_upstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_8_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_8_upstream_byteaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_8_upstream_byteenable : OUT STD_LOGIC;
                 signal niosII_system_burst_8_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_8_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_8_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_8_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_8_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_8_upstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity niosII_system_burst_8_upstream_arbitrator;


architecture europa of niosII_system_burst_8_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_8_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_8_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_8_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_8_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_8_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_8_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_8_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_8_upstream_write :  STD_LOGIC;
                signal module_input120 :  STD_LOGIC;
                signal module_input121 :  STD_LOGIC;
                signal module_input122 :  STD_LOGIC;
                signal module_input123 :  STD_LOGIC;
                signal module_input124 :  STD_LOGIC;
                signal module_input125 :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_8_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_8_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_8_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_8_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_8_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_8_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_8_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_8_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_8_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_8_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_8_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_8_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_8_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_8_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_8_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_8_upstream);
  --assign niosII_system_burst_8_upstream_readdatavalid_from_sa = niosII_system_burst_8_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_8_upstream_readdatavalid_from_sa <= niosII_system_burst_8_upstream_readdatavalid;
  --assign niosII_system_burst_8_upstream_readdata_from_sa = niosII_system_burst_8_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_8_upstream_readdata_from_sa <= niosII_system_burst_8_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_8_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1100100001001000010010000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_8_upstream_waitrequest_from_sa = niosII_system_burst_8_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_8_upstream_waitrequest_from_sa <= niosII_system_burst_8_upstream_waitrequest;
  --niosII_system_burst_8_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_8_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_8_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_8_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_8_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_8_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_8_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_8_upstream;
  --niosII_system_burst_8_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_8_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_8_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_8_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_8_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_8_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_8_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_8_upstream_allgrants <= niosII_system_burst_8_upstream_grant_vector;
  --niosII_system_burst_8_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_8_upstream_end_xfer <= NOT ((niosII_system_burst_8_upstream_waits_for_read OR niosII_system_burst_8_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_8_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_8_upstream <= niosII_system_burst_8_upstream_end_xfer AND (((NOT niosII_system_burst_8_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_8_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_8_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_8_upstream AND niosII_system_burst_8_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_8_upstream AND NOT niosII_system_burst_8_upstream_non_bursting_master_requests));
  --niosII_system_burst_8_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_8_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_8_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_8_upstream_arb_share_counter <= niosII_system_burst_8_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_8_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_8_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_8_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_8_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_8_upstream AND NOT niosII_system_burst_8_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_8_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_8_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_8/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_8_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_8_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_8_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_8_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_8/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_8_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_8_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_8_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_8_upstream <= internal_cpu_data_master_requests_niosII_system_burst_8_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register)))));
  --unique name for niosII_system_burst_8_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_8_upstream_move_on_to_next_transaction <= niosII_system_burst_8_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_8_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_8_upstream, which is an e_mux
  niosII_system_burst_8_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_8_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_8_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_8_upstream : burstcount_fifo_for_niosII_system_burst_8_upstream_module
    port map(
      data_out => niosII_system_burst_8_upstream_transaction_burst_count,
      empty => niosII_system_burst_8_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input120,
      clk => clk,
      data_in => niosII_system_burst_8_upstream_selected_burstcount,
      read => niosII_system_burst_8_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input121,
      write => module_input122
    );

  module_input120 <= std_logic'('0');
  module_input121 <= std_logic'('0');
  module_input122 <= ((in_a_read_cycle AND NOT niosII_system_burst_8_upstream_waits_for_read) AND niosII_system_burst_8_upstream_load_fifo) AND NOT ((niosII_system_burst_8_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_8_upstream_burstcount_fifo_empty));

  --niosII_system_burst_8_upstream current burst minus one, which is an e_assign
  niosII_system_burst_8_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_8_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_8_upstream, which is an e_mux
  niosII_system_burst_8_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_8_upstream_waits_for_read)) AND NOT niosII_system_burst_8_upstream_load_fifo))) = '1'), niosII_system_burst_8_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_8_upstream_waits_for_read) AND niosII_system_burst_8_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_8_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_8_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_8_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_8_upstream_transaction_burst_count, niosII_system_burst_8_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_8_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_8_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_8_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_8_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_8_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_8_upstream_current_burst <= niosII_system_burst_8_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_8_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_8_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_8_upstream_waits_for_read)) AND niosII_system_burst_8_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_8_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_8_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_8_upstream_waits_for_read)) AND NOT niosII_system_burst_8_upstream_load_fifo) OR niosII_system_burst_8_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_8_upstream_load_fifo <= p0_niosII_system_burst_8_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_8_upstream, which is an e_assign
  niosII_system_burst_8_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_8_upstream_current_burst_minus_one)) AND niosII_system_burst_8_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_8_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_8_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_8_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_8_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_8_upstream,
      full => open,
      clear_fifo => module_input123,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_8_upstream,
      read => niosII_system_burst_8_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input124,
      write => module_input125
    );

  module_input123 <= std_logic'('0');
  module_input124 <= std_logic'('0');
  module_input125 <= in_a_read_cycle AND NOT niosII_system_burst_8_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_8_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_8_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_8_upstream <= niosII_system_burst_8_upstream_readdatavalid_from_sa;
  --niosII_system_burst_8_upstream_writedata mux, which is an e_mux
  niosII_system_burst_8_upstream_writedata <= cpu_data_master_writedata (7 DOWNTO 0);
  --byteaddress mux for niosII_system_burst_8/upstream, which is an e_mux
  niosII_system_burst_8_upstream_byteaddress <= cpu_data_master_address_to_slave (1 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_8_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_8_upstream;
  --cpu/data_master saved-grant niosII_system_burst_8/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_8_upstream <= internal_cpu_data_master_requests_niosII_system_burst_8_upstream;
  --allow new arb cycle for niosII_system_burst_8/upstream, which is an e_assign
  niosII_system_burst_8_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_8_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_8_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_8_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_8_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_8_upstream_begins_xfer) = '1'), niosII_system_burst_8_upstream_unreg_firsttransfer, niosII_system_burst_8_upstream_reg_firsttransfer);
  --niosII_system_burst_8_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_8_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_8_upstream_slavearbiterlockenable AND niosII_system_burst_8_upstream_any_continuerequest));
  --niosII_system_burst_8_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_8_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_8_upstream_begins_xfer) = '1' then 
        niosII_system_burst_8_upstream_reg_firsttransfer <= niosII_system_burst_8_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_8_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_8_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_8_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_8_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_8_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_8_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_8_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_8_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_8_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_8_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_8_upstream_begins_xfer) = '1' then 
        niosII_system_burst_8_upstream_bbt_burstcounter <= niosII_system_burst_8_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_8_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_8_upstream_beginbursttransfer_internal <= niosII_system_burst_8_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_8_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_8_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_8_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_8_upstream AND cpu_data_master_read;
  --niosII_system_burst_8_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_8_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_8_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_8_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_8_upstream_address mux, which is an e_mux
  niosII_system_burst_8_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_8_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_niosII_system_burst_8_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_8_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_8_upstream_end_xfer <= niosII_system_burst_8_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_8_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_8_upstream_waits_for_read <= niosII_system_burst_8_upstream_in_a_read_cycle AND internal_niosII_system_burst_8_upstream_waitrequest_from_sa;
  --niosII_system_burst_8_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_8_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_8_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_8_upstream_in_a_read_cycle;
  --niosII_system_burst_8_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_8_upstream_waits_for_write <= niosII_system_burst_8_upstream_in_a_write_cycle AND internal_niosII_system_burst_8_upstream_waitrequest_from_sa;
  --niosII_system_burst_8_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_8_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_8_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_8_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_8_upstream_counter <= std_logic'('0');
  --niosII_system_burst_8_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_8_upstream_byteenable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_8_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_8_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_8_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_8_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_8_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_8_upstream <= internal_cpu_data_master_granted_niosII_system_burst_8_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_8_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_8_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_8_upstream <= internal_cpu_data_master_requests_niosII_system_burst_8_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_8_upstream_burstcount <= internal_niosII_system_burst_8_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_8_upstream_read <= internal_niosII_system_burst_8_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_8_upstream_waitrequest_from_sa <= internal_niosII_system_burst_8_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_8_upstream_write <= internal_niosII_system_burst_8_upstream_write;
--synthesis translate_off
    --niosII_system_burst_8/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line171 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_8_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line171, now);
          write(write_line171, string'(": "));
          write(write_line171, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_8/upstream"));
          write(output, write_line171.all);
          deallocate (write_line171);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_8_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_led_pio_s1_end_xfer : IN STD_LOGIC;
                 signal led_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_8_downstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_8_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_byteenable : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_granted_led_pio_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_qualified_request_led_pio_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_read_data_valid_led_pio_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_requests_led_pio_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_8_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_burst_8_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_8_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_8_downstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_8_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_8_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_8_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_8_downstream_arbitrator;


architecture europa of niosII_system_burst_8_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_8_downstream_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_niosII_system_burst_8_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_8_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_byteenable_last_time :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pre_flush_niosII_system_burst_8_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_8_downstream_qualified_request_led_pio_s1 OR NOT niosII_system_burst_8_downstream_requests_led_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_8_downstream_qualified_request_led_pio_s1 OR NOT niosII_system_burst_8_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_led_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_8_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_8_downstream_qualified_request_led_pio_s1 OR NOT niosII_system_burst_8_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_8_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_8_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_8_downstream_address_to_slave <= niosII_system_burst_8_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_8_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_8_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_8_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_8_downstream_read_data_valid_led_pio_s1)))));
  --niosII_system_burst_8/downstream readdata mux, which is an e_mux
  niosII_system_burst_8_downstream_readdata <= led_pio_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_8_downstream_waitrequest <= NOT niosII_system_burst_8_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_8_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_8_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_8_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_8_downstream_address_to_slave <= internal_niosII_system_burst_8_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_8_downstream_waitrequest <= internal_niosII_system_burst_8_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_8_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_8_downstream_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_8_downstream_address_last_time <= niosII_system_burst_8_downstream_address;
      end if;

    end process;

    --niosII_system_burst_8/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_8_downstream_waitrequest AND ((niosII_system_burst_8_downstream_read OR niosII_system_burst_8_downstream_write));
      end if;

    end process;

    --niosII_system_burst_8_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line172 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_8_downstream_address /= niosII_system_burst_8_downstream_address_last_time))))) = '1' then 
          write(write_line172, now);
          write(write_line172, string'(": "));
          write(write_line172, string'("niosII_system_burst_8_downstream_address did not heed wait!!!"));
          write(output, write_line172.all);
          deallocate (write_line172);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_8_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_8_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_8_downstream_burstcount_last_time <= niosII_system_burst_8_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_8_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line173 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_8_downstream_burstcount) /= std_logic'(niosII_system_burst_8_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line173, now);
          write(write_line173, string'(": "));
          write(write_line173, string'("niosII_system_burst_8_downstream_burstcount did not heed wait!!!"));
          write(output, write_line173.all);
          deallocate (write_line173);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_8_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_8_downstream_byteenable_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_8_downstream_byteenable_last_time <= niosII_system_burst_8_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_8_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line174 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_8_downstream_byteenable) /= std_logic'(niosII_system_burst_8_downstream_byteenable_last_time)))))) = '1' then 
          write(write_line174, now);
          write(write_line174, string'(": "));
          write(write_line174, string'("niosII_system_burst_8_downstream_byteenable did not heed wait!!!"));
          write(output, write_line174.all);
          deallocate (write_line174);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_8_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_8_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_8_downstream_read_last_time <= niosII_system_burst_8_downstream_read;
      end if;

    end process;

    --niosII_system_burst_8_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line175 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_8_downstream_read) /= std_logic'(niosII_system_burst_8_downstream_read_last_time)))))) = '1' then 
          write(write_line175, now);
          write(write_line175, string'(": "));
          write(write_line175, string'("niosII_system_burst_8_downstream_read did not heed wait!!!"));
          write(output, write_line175.all);
          deallocate (write_line175);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_8_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_8_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_8_downstream_write_last_time <= niosII_system_burst_8_downstream_write;
      end if;

    end process;

    --niosII_system_burst_8_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line176 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_8_downstream_write) /= std_logic'(niosII_system_burst_8_downstream_write_last_time)))))) = '1' then 
          write(write_line176, now);
          write(write_line176, string'(": "));
          write(write_line176, string'("niosII_system_burst_8_downstream_write did not heed wait!!!"));
          write(output, write_line176.all);
          deallocate (write_line176);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_8_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_8_downstream_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_8_downstream_writedata_last_time <= niosII_system_burst_8_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_8_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line177 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_8_downstream_writedata /= niosII_system_burst_8_downstream_writedata_last_time)))) AND niosII_system_burst_8_downstream_write)) = '1' then 
          write(write_line177, now);
          write(write_line177, string'(": "));
          write(write_line177, string'("niosII_system_burst_8_downstream_writedata did not heed wait!!!"));
          write(output, write_line177.all);
          deallocate (write_line177);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_niosII_system_burst_9_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_niosII_system_burst_9_upstream_module;


architecture europa of burstcount_fifo_for_niosII_system_burst_9_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_9_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_niosII_system_burst_9_upstream_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_niosII_system_burst_9_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_9_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_burst_9_upstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_9_upstream_readdatavalid : IN STD_LOGIC;
                 signal niosII_system_burst_9_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_niosII_system_burst_9_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_niosII_system_burst_9_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_niosII_system_burst_9_upstream : OUT STD_LOGIC;
                 signal d1_niosII_system_burst_9_upstream_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_9_upstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_9_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_9_upstream_byteaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_9_upstream_byteenable : OUT STD_LOGIC;
                 signal niosII_system_burst_9_upstream_debugaccess : OUT STD_LOGIC;
                 signal niosII_system_burst_9_upstream_read : OUT STD_LOGIC;
                 signal niosII_system_burst_9_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_9_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_burst_9_upstream_write : OUT STD_LOGIC;
                 signal niosII_system_burst_9_upstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity niosII_system_burst_9_upstream_arbitrator;


architecture europa of niosII_system_burst_9_upstream_arbitrator is
component burstcount_fifo_for_niosII_system_burst_9_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_niosII_system_burst_9_upstream_module;

component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_9_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_niosII_system_burst_9_upstream_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal cpu_data_master_saved_grant_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal internal_cpu_data_master_requests_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal internal_niosII_system_burst_9_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_burst_9_upstream_read :  STD_LOGIC;
                signal internal_niosII_system_burst_9_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_system_burst_9_upstream_write :  STD_LOGIC;
                signal module_input126 :  STD_LOGIC;
                signal module_input127 :  STD_LOGIC;
                signal module_input128 :  STD_LOGIC;
                signal module_input129 :  STD_LOGIC;
                signal module_input130 :  STD_LOGIC;
                signal module_input131 :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_allgrants :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_any_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_arb_share_counter :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_9_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_9_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_9_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_9_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_begins_xfer :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_9_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_9_upstream_end_xfer :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_grant_vector :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_load_fifo :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_9_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_9_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_9_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_9_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_waits_for_read :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_waits_for_write :  STD_LOGIC;
                signal p0_niosII_system_burst_9_upstream_load_fifo :  STD_LOGIC;
                signal shifted_address_to_niosII_system_burst_9_upstream_from_cpu_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_niosII_system_burst_9_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_burst_9_upstream_end_xfer;
    end if;

  end process;

  niosII_system_burst_9_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_niosII_system_burst_9_upstream);
  --assign niosII_system_burst_9_upstream_readdatavalid_from_sa = niosII_system_burst_9_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_9_upstream_readdatavalid_from_sa <= niosII_system_burst_9_upstream_readdatavalid;
  --assign niosII_system_burst_9_upstream_readdata_from_sa = niosII_system_burst_9_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_burst_9_upstream_readdata_from_sa <= niosII_system_burst_9_upstream_readdata;
  internal_cpu_data_master_requests_niosII_system_burst_9_upstream <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1100100001001000010100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign niosII_system_burst_9_upstream_waitrequest_from_sa = niosII_system_burst_9_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_burst_9_upstream_waitrequest_from_sa <= niosII_system_burst_9_upstream_waitrequest;
  --niosII_system_burst_9_upstream_arb_share_counter set values, which is an e_mux
  niosII_system_burst_9_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_9_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((cpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 8);
  --niosII_system_burst_9_upstream_non_bursting_master_requests mux, which is an e_mux
  niosII_system_burst_9_upstream_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_burst_9_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_burst_9_upstream_any_bursting_master_saved_grant <= cpu_data_master_saved_grant_niosII_system_burst_9_upstream;
  --niosII_system_burst_9_upstream_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_burst_9_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_burst_9_upstream_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_9_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_burst_9_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000") & (niosII_system_burst_9_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 8);
  --niosII_system_burst_9_upstream_allgrants all slave grants, which is an e_mux
  niosII_system_burst_9_upstream_allgrants <= niosII_system_burst_9_upstream_grant_vector;
  --niosII_system_burst_9_upstream_end_xfer assignment, which is an e_assign
  niosII_system_burst_9_upstream_end_xfer <= NOT ((niosII_system_burst_9_upstream_waits_for_read OR niosII_system_burst_9_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_burst_9_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_burst_9_upstream <= niosII_system_burst_9_upstream_end_xfer AND (((NOT niosII_system_burst_9_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_burst_9_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_burst_9_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_burst_9_upstream AND niosII_system_burst_9_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_9_upstream AND NOT niosII_system_burst_9_upstream_non_bursting_master_requests));
  --niosII_system_burst_9_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_9_upstream_arb_share_counter <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_9_upstream_arb_counter_enable) = '1' then 
        niosII_system_burst_9_upstream_arb_share_counter <= niosII_system_burst_9_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_burst_9_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_9_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_burst_9_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_burst_9_upstream)) OR ((end_xfer_arb_share_counter_term_niosII_system_burst_9_upstream AND NOT niosII_system_burst_9_upstream_non_bursting_master_requests)))) = '1' then 
        niosII_system_burst_9_upstream_slavearbiterlockenable <= or_reduce(niosII_system_burst_9_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master niosII_system_burst_9/upstream arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= niosII_system_burst_9_upstream_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --niosII_system_burst_9_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_burst_9_upstream_slavearbiterlockenable2 <= or_reduce(niosII_system_burst_9_upstream_arb_share_counter_next_value);
  --cpu/data_master niosII_system_burst_9/upstream arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= niosII_system_burst_9_upstream_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --niosII_system_burst_9_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_burst_9_upstream_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_niosII_system_burst_9_upstream <= internal_cpu_data_master_requests_niosII_system_burst_9_upstream AND NOT ((cpu_data_master_read AND (((((((((((((((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_latency_counter))))))) OR (cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register)) OR (cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register)))));
  --unique name for niosII_system_burst_9_upstream_move_on_to_next_transaction, which is an e_assign
  niosII_system_burst_9_upstream_move_on_to_next_transaction <= niosII_system_burst_9_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_9_upstream_load_fifo;
  --the currently selected burstcount for niosII_system_burst_9_upstream, which is an e_mux
  niosII_system_burst_9_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_9_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_niosII_system_burst_9_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_niosII_system_burst_9_upstream : burstcount_fifo_for_niosII_system_burst_9_upstream_module
    port map(
      data_out => niosII_system_burst_9_upstream_transaction_burst_count,
      empty => niosII_system_burst_9_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input126,
      clk => clk,
      data_in => niosII_system_burst_9_upstream_selected_burstcount,
      read => niosII_system_burst_9_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input127,
      write => module_input128
    );

  module_input126 <= std_logic'('0');
  module_input127 <= std_logic'('0');
  module_input128 <= ((in_a_read_cycle AND NOT niosII_system_burst_9_upstream_waits_for_read) AND niosII_system_burst_9_upstream_load_fifo) AND NOT ((niosII_system_burst_9_upstream_this_cycle_is_the_last_burst AND niosII_system_burst_9_upstream_burstcount_fifo_empty));

  --niosII_system_burst_9_upstream current burst minus one, which is an e_assign
  niosII_system_burst_9_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_9_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for niosII_system_burst_9_upstream, which is an e_mux
  niosII_system_burst_9_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_9_upstream_waits_for_read)) AND NOT niosII_system_burst_9_upstream_load_fifo))) = '1'), niosII_system_burst_9_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_9_upstream_waits_for_read) AND niosII_system_burst_9_upstream_this_cycle_is_the_last_burst) AND niosII_system_burst_9_upstream_burstcount_fifo_empty))) = '1'), niosII_system_burst_9_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((niosII_system_burst_9_upstream_this_cycle_is_the_last_burst)) = '1'), niosII_system_burst_9_upstream_transaction_burst_count, niosII_system_burst_9_upstream_current_burst_minus_one)));
  --the current burst count for niosII_system_burst_9_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_9_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((niosII_system_burst_9_upstream_readdatavalid_from_sa OR ((NOT niosII_system_burst_9_upstream_load_fifo AND ((in_a_read_cycle AND NOT niosII_system_burst_9_upstream_waits_for_read)))))) = '1' then 
        niosII_system_burst_9_upstream_current_burst <= niosII_system_burst_9_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_niosII_system_burst_9_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT niosII_system_burst_9_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_9_upstream_waits_for_read)) AND niosII_system_burst_9_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_system_burst_9_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_9_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT niosII_system_burst_9_upstream_waits_for_read)) AND NOT niosII_system_burst_9_upstream_load_fifo) OR niosII_system_burst_9_upstream_this_cycle_is_the_last_burst)) = '1' then 
        niosII_system_burst_9_upstream_load_fifo <= p0_niosII_system_burst_9_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for niosII_system_burst_9_upstream, which is an e_assign
  niosII_system_burst_9_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(niosII_system_burst_9_upstream_current_burst_minus_one)) AND niosII_system_burst_9_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_niosII_system_burst_9_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_niosII_system_burst_9_upstream : rdv_fifo_for_cpu_data_master_to_niosII_system_burst_9_upstream_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_niosII_system_burst_9_upstream,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_niosII_system_burst_9_upstream,
      full => open,
      clear_fifo => module_input129,
      clk => clk,
      data_in => internal_cpu_data_master_granted_niosII_system_burst_9_upstream,
      read => niosII_system_burst_9_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input130,
      write => module_input131
    );

  module_input129 <= std_logic'('0');
  module_input130 <= std_logic'('0');
  module_input131 <= in_a_read_cycle AND NOT niosII_system_burst_9_upstream_waits_for_read;

  cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register <= NOT cpu_data_master_rdv_fifo_empty_niosII_system_burst_9_upstream;
  --local readdatavalid cpu_data_master_read_data_valid_niosII_system_burst_9_upstream, which is an e_mux
  cpu_data_master_read_data_valid_niosII_system_burst_9_upstream <= niosII_system_burst_9_upstream_readdatavalid_from_sa;
  --niosII_system_burst_9_upstream_writedata mux, which is an e_mux
  niosII_system_burst_9_upstream_writedata <= cpu_data_master_writedata (7 DOWNTO 0);
  --byteaddress mux for niosII_system_burst_9/upstream, which is an e_mux
  niosII_system_burst_9_upstream_byteaddress <= cpu_data_master_address_to_slave (1 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_niosII_system_burst_9_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_9_upstream;
  --cpu/data_master saved-grant niosII_system_burst_9/upstream, which is an e_assign
  cpu_data_master_saved_grant_niosII_system_burst_9_upstream <= internal_cpu_data_master_requests_niosII_system_burst_9_upstream;
  --allow new arb cycle for niosII_system_burst_9/upstream, which is an e_assign
  niosII_system_burst_9_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_burst_9_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_burst_9_upstream_master_qreq_vector <= std_logic'('1');
  --niosII_system_burst_9_upstream_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_9_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_burst_9_upstream_begins_xfer) = '1'), niosII_system_burst_9_upstream_unreg_firsttransfer, niosII_system_burst_9_upstream_reg_firsttransfer);
  --niosII_system_burst_9_upstream_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_burst_9_upstream_unreg_firsttransfer <= NOT ((niosII_system_burst_9_upstream_slavearbiterlockenable AND niosII_system_burst_9_upstream_any_continuerequest));
  --niosII_system_burst_9_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_9_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_9_upstream_begins_xfer) = '1' then 
        niosII_system_burst_9_upstream_reg_firsttransfer <= niosII_system_burst_9_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_burst_9_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  niosII_system_burst_9_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_9_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_9_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_niosII_system_burst_9_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_niosII_system_burst_9_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_9_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_9_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --niosII_system_burst_9_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_9_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_burst_9_upstream_begins_xfer) = '1' then 
        niosII_system_burst_9_upstream_bbt_burstcounter <= niosII_system_burst_9_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --niosII_system_burst_9_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_burst_9_upstream_beginbursttransfer_internal <= niosII_system_burst_9_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (niosII_system_burst_9_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --niosII_system_burst_9_upstream_read assignment, which is an e_mux
  internal_niosII_system_burst_9_upstream_read <= internal_cpu_data_master_granted_niosII_system_burst_9_upstream AND cpu_data_master_read;
  --niosII_system_burst_9_upstream_write assignment, which is an e_mux
  internal_niosII_system_burst_9_upstream_write <= internal_cpu_data_master_granted_niosII_system_burst_9_upstream AND cpu_data_master_write;
  shifted_address_to_niosII_system_burst_9_upstream_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --niosII_system_burst_9_upstream_address mux, which is an e_mux
  niosII_system_burst_9_upstream_address <= A_EXT (A_SRL(shifted_address_to_niosII_system_burst_9_upstream_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_niosII_system_burst_9_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_burst_9_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_burst_9_upstream_end_xfer <= niosII_system_burst_9_upstream_end_xfer;
    end if;

  end process;

  --niosII_system_burst_9_upstream_waits_for_read in a cycle, which is an e_mux
  niosII_system_burst_9_upstream_waits_for_read <= niosII_system_burst_9_upstream_in_a_read_cycle AND internal_niosII_system_burst_9_upstream_waitrequest_from_sa;
  --niosII_system_burst_9_upstream_in_a_read_cycle assignment, which is an e_assign
  niosII_system_burst_9_upstream_in_a_read_cycle <= internal_cpu_data_master_granted_niosII_system_burst_9_upstream AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_burst_9_upstream_in_a_read_cycle;
  --niosII_system_burst_9_upstream_waits_for_write in a cycle, which is an e_mux
  niosII_system_burst_9_upstream_waits_for_write <= niosII_system_burst_9_upstream_in_a_write_cycle AND internal_niosII_system_burst_9_upstream_waitrequest_from_sa;
  --niosII_system_burst_9_upstream_in_a_write_cycle assignment, which is an e_assign
  niosII_system_burst_9_upstream_in_a_write_cycle <= internal_cpu_data_master_granted_niosII_system_burst_9_upstream AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_burst_9_upstream_in_a_write_cycle;
  wait_for_niosII_system_burst_9_upstream_counter <= std_logic'('0');
  --niosII_system_burst_9_upstream_byteenable byte enable port mux, which is an e_mux
  niosII_system_burst_9_upstream_byteenable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_9_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --burstcount mux, which is an e_mux
  internal_niosII_system_burst_9_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_9_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  niosII_system_burst_9_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_niosII_system_burst_9_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_niosII_system_burst_9_upstream <= internal_cpu_data_master_granted_niosII_system_burst_9_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_niosII_system_burst_9_upstream <= internal_cpu_data_master_qualified_request_niosII_system_burst_9_upstream;
  --vhdl renameroo for output signals
  cpu_data_master_requests_niosII_system_burst_9_upstream <= internal_cpu_data_master_requests_niosII_system_burst_9_upstream;
  --vhdl renameroo for output signals
  niosII_system_burst_9_upstream_burstcount <= internal_niosII_system_burst_9_upstream_burstcount;
  --vhdl renameroo for output signals
  niosII_system_burst_9_upstream_read <= internal_niosII_system_burst_9_upstream_read;
  --vhdl renameroo for output signals
  niosII_system_burst_9_upstream_waitrequest_from_sa <= internal_niosII_system_burst_9_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_system_burst_9_upstream_write <= internal_niosII_system_burst_9_upstream_write;
--synthesis translate_off
    --niosII_system_burst_9/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --cpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line178 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_cpu_data_master_requests_niosII_system_burst_9_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line178, now);
          write(write_line178, string'(": "));
          write(write_line178, string'("cpu/data_master drove 0 on its 'burstcount' port while accessing slave niosII_system_burst_9/upstream"));
          write(output, write_line178.all);
          deallocate (write_line178);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_burst_9_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_switch_s1_end_xfer : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_9_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_byteenable : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_granted_switch_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_qualified_request_switch_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_read_data_valid_switch_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_requests_switch_s1 : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal switch_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- outputs:
                 signal niosII_system_burst_9_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_9_downstream_latency_counter : OUT STD_LOGIC;
                 signal niosII_system_burst_9_downstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_9_downstream_readdatavalid : OUT STD_LOGIC;
                 signal niosII_system_burst_9_downstream_reset_n : OUT STD_LOGIC;
                 signal niosII_system_burst_9_downstream_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_burst_9_downstream_arbitrator;


architecture europa of niosII_system_burst_9_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_burst_9_downstream_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_niosII_system_burst_9_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_9_downstream_burstcount_last_time :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_byteenable_last_time :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_read_last_time :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_run :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_write_last_time :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pre_flush_niosII_system_burst_9_downstream_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_9_downstream_qualified_request_switch_s1 OR NOT niosII_system_burst_9_downstream_requests_switch_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_9_downstream_qualified_request_switch_s1 OR NOT niosII_system_burst_9_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_switch_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_9_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_burst_9_downstream_qualified_request_switch_s1 OR NOT niosII_system_burst_9_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_9_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_burst_9_downstream_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_burst_9_downstream_address_to_slave <= niosII_system_burst_9_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_niosII_system_burst_9_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  niosII_system_burst_9_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_niosII_system_burst_9_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_9_downstream_read_data_valid_switch_s1)))));
  --niosII_system_burst_9/downstream readdata mux, which is an e_mux
  niosII_system_burst_9_downstream_readdata <= switch_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_burst_9_downstream_waitrequest <= NOT niosII_system_burst_9_downstream_run;
  --latent max counter, which is an e_assign
  niosII_system_burst_9_downstream_latency_counter <= std_logic'('0');
  --niosII_system_burst_9_downstream_reset_n assignment, which is an e_assign
  niosII_system_burst_9_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_burst_9_downstream_address_to_slave <= internal_niosII_system_burst_9_downstream_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_9_downstream_waitrequest <= internal_niosII_system_burst_9_downstream_waitrequest;
--synthesis translate_off
    --niosII_system_burst_9_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_9_downstream_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_system_burst_9_downstream_address_last_time <= niosII_system_burst_9_downstream_address;
      end if;

    end process;

    --niosII_system_burst_9/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_burst_9_downstream_waitrequest AND ((niosII_system_burst_9_downstream_read OR niosII_system_burst_9_downstream_write));
      end if;

    end process;

    --niosII_system_burst_9_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line179 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_9_downstream_address /= niosII_system_burst_9_downstream_address_last_time))))) = '1' then 
          write(write_line179, now);
          write(write_line179, string'(": "));
          write(write_line179, string'("niosII_system_burst_9_downstream_address did not heed wait!!!"));
          write(output, write_line179.all);
          deallocate (write_line179);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_9_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_9_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_9_downstream_burstcount_last_time <= niosII_system_burst_9_downstream_burstcount;
      end if;

    end process;

    --niosII_system_burst_9_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line180 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_9_downstream_burstcount) /= std_logic'(niosII_system_burst_9_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line180, now);
          write(write_line180, string'(": "));
          write(write_line180, string'("niosII_system_burst_9_downstream_burstcount did not heed wait!!!"));
          write(output, write_line180.all);
          deallocate (write_line180);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_9_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_9_downstream_byteenable_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_9_downstream_byteenable_last_time <= niosII_system_burst_9_downstream_byteenable;
      end if;

    end process;

    --niosII_system_burst_9_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line181 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_9_downstream_byteenable) /= std_logic'(niosII_system_burst_9_downstream_byteenable_last_time)))))) = '1' then 
          write(write_line181, now);
          write(write_line181, string'(": "));
          write(write_line181, string'("niosII_system_burst_9_downstream_byteenable did not heed wait!!!"));
          write(output, write_line181.all);
          deallocate (write_line181);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_9_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_9_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_9_downstream_read_last_time <= niosII_system_burst_9_downstream_read;
      end if;

    end process;

    --niosII_system_burst_9_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line182 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_9_downstream_read) /= std_logic'(niosII_system_burst_9_downstream_read_last_time)))))) = '1' then 
          write(write_line182, now);
          write(write_line182, string'(": "));
          write(write_line182, string'("niosII_system_burst_9_downstream_read did not heed wait!!!"));
          write(output, write_line182.all);
          deallocate (write_line182);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_9_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_9_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_burst_9_downstream_write_last_time <= niosII_system_burst_9_downstream_write;
      end if;

    end process;

    --niosII_system_burst_9_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line183 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_burst_9_downstream_write) /= std_logic'(niosII_system_burst_9_downstream_write_last_time)))))) = '1' then 
          write(write_line183, now);
          write(write_line183, string'(": "));
          write(write_line183, string'("niosII_system_burst_9_downstream_write did not heed wait!!!"));
          write(output, write_line183.all);
          deallocate (write_line183);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_9_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_burst_9_downstream_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        niosII_system_burst_9_downstream_writedata_last_time <= niosII_system_burst_9_downstream_writedata;
      end if;

    end process;

    --niosII_system_burst_9_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line184 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_burst_9_downstream_writedata /= niosII_system_burst_9_downstream_writedata_last_time)))) AND niosII_system_burst_9_downstream_write)) = '1' then 
          write(write_line184, now);
          write(write_line184, string'(": "));
          write(write_line184, string'("niosII_system_burst_9_downstream_writedata did not heed wait!!!"));
          write(output, write_line184.all);
          deallocate (write_line184);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_clock_0_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_21_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_21_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_21_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_21_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_21_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_clock_0_in_endofpacket : IN STD_LOGIC;
                 signal niosII_system_clock_0_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_clock_0_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_niosII_system_clock_0_in_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in : OUT STD_LOGIC;
                 signal niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in : OUT STD_LOGIC;
                 signal niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in : OUT STD_LOGIC;
                 signal niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in : OUT STD_LOGIC;
                 signal niosII_system_clock_0_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal niosII_system_clock_0_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_clock_0_in_read : OUT STD_LOGIC;
                 signal niosII_system_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_clock_0_in_reset_n : OUT STD_LOGIC;
                 signal niosII_system_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_system_clock_0_in_write : OUT STD_LOGIC;
                 signal niosII_system_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity niosII_system_clock_0_in_arbitrator;


architecture europa of niosII_system_clock_0_in_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_system_clock_0_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in :  STD_LOGIC;
                signal internal_niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in :  STD_LOGIC;
                signal internal_niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in :  STD_LOGIC;
                signal internal_niosII_system_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_saved_grant_niosII_system_clock_0_in :  STD_LOGIC;
                signal niosII_system_clock_0_in_allgrants :  STD_LOGIC;
                signal niosII_system_clock_0_in_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_system_clock_0_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_system_clock_0_in_any_continuerequest :  STD_LOGIC;
                signal niosII_system_clock_0_in_arb_counter_enable :  STD_LOGIC;
                signal niosII_system_clock_0_in_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_clock_0_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_clock_0_in_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_clock_0_in_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_system_clock_0_in_begins_xfer :  STD_LOGIC;
                signal niosII_system_clock_0_in_end_xfer :  STD_LOGIC;
                signal niosII_system_clock_0_in_firsttransfer :  STD_LOGIC;
                signal niosII_system_clock_0_in_grant_vector :  STD_LOGIC;
                signal niosII_system_clock_0_in_in_a_read_cycle :  STD_LOGIC;
                signal niosII_system_clock_0_in_in_a_write_cycle :  STD_LOGIC;
                signal niosII_system_clock_0_in_master_qreq_vector :  STD_LOGIC;
                signal niosII_system_clock_0_in_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_system_clock_0_in_reg_firsttransfer :  STD_LOGIC;
                signal niosII_system_clock_0_in_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_system_clock_0_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_system_clock_0_in_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_system_clock_0_in_waits_for_read :  STD_LOGIC;
                signal niosII_system_clock_0_in_waits_for_write :  STD_LOGIC;
                signal wait_for_niosII_system_clock_0_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_system_clock_0_in_end_xfer;
    end if;

  end process;

  niosII_system_clock_0_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in);
  --assign niosII_system_clock_0_in_readdata_from_sa = niosII_system_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_clock_0_in_readdata_from_sa <= niosII_system_clock_0_in_readdata;
  internal_niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_21_downstream_read OR niosII_system_burst_21_downstream_write)))))));
  --assign niosII_system_clock_0_in_waitrequest_from_sa = niosII_system_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_system_clock_0_in_waitrequest_from_sa <= niosII_system_clock_0_in_waitrequest;
  --niosII_system_clock_0_in_arb_share_counter set values, which is an e_mux
  niosII_system_clock_0_in_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_21_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --niosII_system_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  niosII_system_clock_0_in_non_bursting_master_requests <= std_logic'('0');
  --niosII_system_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_system_clock_0_in_any_bursting_master_saved_grant <= niosII_system_burst_21_downstream_saved_grant_niosII_system_clock_0_in;
  --niosII_system_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  niosII_system_clock_0_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_system_clock_0_in_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_clock_0_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_system_clock_0_in_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (niosII_system_clock_0_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --niosII_system_clock_0_in_allgrants all slave grants, which is an e_mux
  niosII_system_clock_0_in_allgrants <= niosII_system_clock_0_in_grant_vector;
  --niosII_system_clock_0_in_end_xfer assignment, which is an e_assign
  niosII_system_clock_0_in_end_xfer <= NOT ((niosII_system_clock_0_in_waits_for_read OR niosII_system_clock_0_in_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_system_clock_0_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_system_clock_0_in <= niosII_system_clock_0_in_end_xfer AND (((NOT niosII_system_clock_0_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_system_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_system_clock_0_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_system_clock_0_in AND niosII_system_clock_0_in_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_system_clock_0_in AND NOT niosII_system_clock_0_in_non_bursting_master_requests));
  --niosII_system_clock_0_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_clock_0_in_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_clock_0_in_arb_counter_enable) = '1' then 
        niosII_system_clock_0_in_arb_share_counter <= niosII_system_clock_0_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_system_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_clock_0_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_system_clock_0_in_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_system_clock_0_in)) OR ((end_xfer_arb_share_counter_term_niosII_system_clock_0_in AND NOT niosII_system_clock_0_in_non_bursting_master_requests)))) = '1' then 
        niosII_system_clock_0_in_slavearbiterlockenable <= or_reduce(niosII_system_clock_0_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_21/downstream niosII_system_clock_0/in arbiterlock, which is an e_assign
  niosII_system_burst_21_downstream_arbiterlock <= niosII_system_clock_0_in_slavearbiterlockenable AND niosII_system_burst_21_downstream_continuerequest;
  --niosII_system_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_system_clock_0_in_slavearbiterlockenable2 <= or_reduce(niosII_system_clock_0_in_arb_share_counter_next_value);
  --niosII_system_burst_21/downstream niosII_system_clock_0/in arbiterlock2, which is an e_assign
  niosII_system_burst_21_downstream_arbiterlock2 <= niosII_system_clock_0_in_slavearbiterlockenable2 AND niosII_system_burst_21_downstream_continuerequest;
  --niosII_system_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_system_clock_0_in_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_21_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_21_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in <= internal_niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in AND NOT ((niosII_system_burst_21_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_21_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in, which is an e_mux
  niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in <= (internal_niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in AND niosII_system_burst_21_downstream_read) AND NOT niosII_system_clock_0_in_waits_for_read;
  --niosII_system_clock_0_in_writedata mux, which is an e_mux
  niosII_system_clock_0_in_writedata <= niosII_system_burst_21_downstream_writedata;
  --assign niosII_system_clock_0_in_endofpacket_from_sa = niosII_system_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_system_clock_0_in_endofpacket_from_sa <= niosII_system_clock_0_in_endofpacket;
  --master is always granted when requested
  internal_niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in <= internal_niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in;
  --niosII_system_burst_21/downstream saved-grant niosII_system_clock_0/in, which is an e_assign
  niosII_system_burst_21_downstream_saved_grant_niosII_system_clock_0_in <= internal_niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in;
  --allow new arb cycle for niosII_system_clock_0/in, which is an e_assign
  niosII_system_clock_0_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_system_clock_0_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_system_clock_0_in_master_qreq_vector <= std_logic'('1');
  --niosII_system_clock_0_in_reset_n assignment, which is an e_assign
  niosII_system_clock_0_in_reset_n <= reset_n;
  --niosII_system_clock_0_in_firsttransfer first transaction, which is an e_assign
  niosII_system_clock_0_in_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_system_clock_0_in_begins_xfer) = '1'), niosII_system_clock_0_in_unreg_firsttransfer, niosII_system_clock_0_in_reg_firsttransfer);
  --niosII_system_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  niosII_system_clock_0_in_unreg_firsttransfer <= NOT ((niosII_system_clock_0_in_slavearbiterlockenable AND niosII_system_clock_0_in_any_continuerequest));
  --niosII_system_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_clock_0_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_system_clock_0_in_begins_xfer) = '1' then 
        niosII_system_clock_0_in_reg_firsttransfer <= niosII_system_clock_0_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_system_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_system_clock_0_in_beginbursttransfer_internal <= niosII_system_clock_0_in_begins_xfer;
  --niosII_system_clock_0_in_read assignment, which is an e_mux
  niosII_system_clock_0_in_read <= internal_niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in AND niosII_system_burst_21_downstream_read;
  --niosII_system_clock_0_in_write assignment, which is an e_mux
  niosII_system_clock_0_in_write <= internal_niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in AND niosII_system_burst_21_downstream_write;
  --niosII_system_clock_0_in_address mux, which is an e_mux
  niosII_system_clock_0_in_address <= niosII_system_burst_21_downstream_address_to_slave;
  --slaveid niosII_system_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  niosII_system_clock_0_in_nativeaddress <= niosII_system_burst_21_downstream_nativeaddress (1 DOWNTO 0);
  --d1_niosII_system_clock_0_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_system_clock_0_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_system_clock_0_in_end_xfer <= niosII_system_clock_0_in_end_xfer;
    end if;

  end process;

  --niosII_system_clock_0_in_waits_for_read in a cycle, which is an e_mux
  niosII_system_clock_0_in_waits_for_read <= niosII_system_clock_0_in_in_a_read_cycle AND internal_niosII_system_clock_0_in_waitrequest_from_sa;
  --niosII_system_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  niosII_system_clock_0_in_in_a_read_cycle <= internal_niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in AND niosII_system_burst_21_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_system_clock_0_in_in_a_read_cycle;
  --niosII_system_clock_0_in_waits_for_write in a cycle, which is an e_mux
  niosII_system_clock_0_in_waits_for_write <= niosII_system_clock_0_in_in_a_write_cycle AND internal_niosII_system_clock_0_in_waitrequest_from_sa;
  --niosII_system_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  niosII_system_clock_0_in_in_a_write_cycle <= internal_niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in AND niosII_system_burst_21_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_system_clock_0_in_in_a_write_cycle;
  wait_for_niosII_system_clock_0_in_counter <= std_logic'('0');
  --niosII_system_clock_0_in_byteenable byte enable port mux, which is an e_mux
  niosII_system_clock_0_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_21_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in <= internal_niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in;
  --vhdl renameroo for output signals
  niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in <= internal_niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in;
  --vhdl renameroo for output signals
  niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in <= internal_niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in;
  --vhdl renameroo for output signals
  niosII_system_clock_0_in_waitrequest_from_sa <= internal_niosII_system_clock_0_in_waitrequest_from_sa;
--synthesis translate_off
    --niosII_system_clock_0/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_21/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line185 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_21_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line185, now);
          write(write_line185, string'(": "));
          write(write_line185, string'("niosII_system_burst_21/downstream drove 0 on its 'arbitrationshare' port while accessing slave niosII_system_clock_0/in"));
          write(output, write_line185.all);
          deallocate (write_line185);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_21/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line186 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_21_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line186, now);
          write(write_line186, string'(": "));
          write(write_line186, string'("niosII_system_burst_21/downstream drove 0 on its 'burstcount' port while accessing slave niosII_system_clock_0/in"));
          write(output, write_line186.all);
          deallocate (write_line186);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_system_clock_0_out_arbitrator is 
        port (
              -- inputs:
                 signal altpll_inst_pll_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_altpll_inst_pll_slave_end_xfer : IN STD_LOGIC;
                 signal niosII_system_clock_0_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_clock_0_out_granted_altpll_inst_pll_slave : IN STD_LOGIC;
                 signal niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave : IN STD_LOGIC;
                 signal niosII_system_clock_0_out_read : IN STD_LOGIC;
                 signal niosII_system_clock_0_out_read_data_valid_altpll_inst_pll_slave : IN STD_LOGIC;
                 signal niosII_system_clock_0_out_requests_altpll_inst_pll_slave : IN STD_LOGIC;
                 signal niosII_system_clock_0_out_write : IN STD_LOGIC;
                 signal niosII_system_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_system_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_system_clock_0_out_reset_n : OUT STD_LOGIC;
                 signal niosII_system_clock_0_out_waitrequest : OUT STD_LOGIC
              );
end entity niosII_system_clock_0_out_arbitrator;


architecture europa of niosII_system_clock_0_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_system_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_system_clock_0_out_waitrequest :  STD_LOGIC;
                signal niosII_system_clock_0_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_clock_0_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_clock_0_out_read_last_time :  STD_LOGIC;
                signal niosII_system_clock_0_out_run :  STD_LOGIC;
                signal niosII_system_clock_0_out_write_last_time :  STD_LOGIC;
                signal niosII_system_clock_0_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave OR NOT ((niosII_system_clock_0_out_read OR niosII_system_clock_0_out_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_clock_0_out_read OR niosII_system_clock_0_out_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave OR NOT ((niosII_system_clock_0_out_read OR niosII_system_clock_0_out_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_clock_0_out_read OR niosII_system_clock_0_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_system_clock_0_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_system_clock_0_out_address_to_slave <= niosII_system_clock_0_out_address;
  --niosII_system_clock_0/out readdata mux, which is an e_mux
  niosII_system_clock_0_out_readdata <= altpll_inst_pll_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_system_clock_0_out_waitrequest <= NOT niosII_system_clock_0_out_run;
  --niosII_system_clock_0_out_reset_n assignment, which is an e_assign
  niosII_system_clock_0_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_system_clock_0_out_address_to_slave <= internal_niosII_system_clock_0_out_address_to_slave;
  --vhdl renameroo for output signals
  niosII_system_clock_0_out_waitrequest <= internal_niosII_system_clock_0_out_waitrequest;
--synthesis translate_off
    --niosII_system_clock_0_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_clock_0_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_clock_0_out_address_last_time <= niosII_system_clock_0_out_address;
      end if;

    end process;

    --niosII_system_clock_0/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_system_clock_0_out_waitrequest AND ((niosII_system_clock_0_out_read OR niosII_system_clock_0_out_write));
      end if;

    end process;

    --niosII_system_clock_0_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line187 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_clock_0_out_address /= niosII_system_clock_0_out_address_last_time))))) = '1' then 
          write(write_line187, now);
          write(write_line187, string'(": "));
          write(write_line187, string'("niosII_system_clock_0_out_address did not heed wait!!!"));
          write(output, write_line187.all);
          deallocate (write_line187);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_clock_0_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_clock_0_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_system_clock_0_out_byteenable_last_time <= niosII_system_clock_0_out_byteenable;
      end if;

    end process;

    --niosII_system_clock_0_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line188 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_system_clock_0_out_byteenable /= niosII_system_clock_0_out_byteenable_last_time))))) = '1' then 
          write(write_line188, now);
          write(write_line188, string'(": "));
          write(write_line188, string'("niosII_system_clock_0_out_byteenable did not heed wait!!!"));
          write(output, write_line188.all);
          deallocate (write_line188);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_clock_0_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_clock_0_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_clock_0_out_read_last_time <= niosII_system_clock_0_out_read;
      end if;

    end process;

    --niosII_system_clock_0_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line189 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_clock_0_out_read) /= std_logic'(niosII_system_clock_0_out_read_last_time)))))) = '1' then 
          write(write_line189, now);
          write(write_line189, string'(": "));
          write(write_line189, string'("niosII_system_clock_0_out_read did not heed wait!!!"));
          write(output, write_line189.all);
          deallocate (write_line189);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_clock_0_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_clock_0_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_system_clock_0_out_write_last_time <= niosII_system_clock_0_out_write;
      end if;

    end process;

    --niosII_system_clock_0_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line190 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_system_clock_0_out_write) /= std_logic'(niosII_system_clock_0_out_write_last_time)))))) = '1' then 
          write(write_line190, now);
          write(write_line190, string'(": "));
          write(write_line190, string'("niosII_system_clock_0_out_write did not heed wait!!!"));
          write(output, write_line190.all);
          deallocate (write_line190);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_clock_0_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_system_clock_0_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_system_clock_0_out_writedata_last_time <= niosII_system_clock_0_out_writedata;
      end if;

    end process;

    --niosII_system_clock_0_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line191 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_system_clock_0_out_writedata /= niosII_system_clock_0_out_writedata_last_time)))) AND niosII_system_clock_0_out_write)) = '1' then 
          write(write_line191, now);
          write(write_line191, string'(": "));
          write(write_line191, string'("niosII_system_clock_0_out_writedata did not heed wait!!!"));
          write(output, write_line191.all);
          deallocate (write_line191);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_niosII_system_burst_10_downstream_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_niosII_system_burst_10_downstream_to_sdram_s1_module;


architecture europa of rdv_fifo_for_niosII_system_burst_10_downstream_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_niosII_system_burst_11_downstream_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_niosII_system_burst_11_downstream_to_sdram_s1_module;


architecture europa of rdv_fifo_for_niosII_system_burst_11_downstream_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sdram_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_address_to_slave : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal niosII_system_burst_10_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_10_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_10_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_10_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_11_downstream_address_to_slave : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal niosII_system_burst_11_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_11_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_11_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_11_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_readdatavalid : IN STD_LOGIC;
                 signal sdram_s1_waitrequest : IN STD_LOGIC;

              -- outputs:
                 signal d1_sdram_s1_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_10_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_10_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_10_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_10_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal niosII_system_burst_10_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_11_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_11_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_11_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_11_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal niosII_system_burst_11_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                 signal sdram_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal sdram_s1_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sdram_s1_chipselect : OUT STD_LOGIC;
                 signal sdram_s1_read_n : OUT STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_reset_n : OUT STD_LOGIC;
                 signal sdram_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal sdram_s1_write_n : OUT STD_LOGIC;
                 signal sdram_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sdram_s1_arbitrator;


architecture europa of sdram_s1_arbitrator is
component rdv_fifo_for_niosII_system_burst_10_downstream_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_niosII_system_burst_10_downstream_to_sdram_s1_module;

component rdv_fifo_for_niosII_system_burst_11_downstream_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_niosII_system_burst_11_downstream_to_sdram_s1_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sdram_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_10_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_10_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_10_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_11_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_11_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_11_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal internal_sdram_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_niosII_system_burst_10_downstream_granted_slave_sdram_s1 :  STD_LOGIC;
                signal last_cycle_niosII_system_burst_11_downstream_granted_slave_sdram_s1 :  STD_LOGIC;
                signal module_input132 :  STD_LOGIC;
                signal module_input133 :  STD_LOGIC;
                signal module_input134 :  STD_LOGIC;
                signal module_input135 :  STD_LOGIC;
                signal module_input136 :  STD_LOGIC;
                signal module_input137 :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_saved_grant_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_saved_grant_sdram_s1 :  STD_LOGIC;
                signal sdram_s1_allgrants :  STD_LOGIC;
                signal sdram_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sdram_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sdram_s1_any_continuerequest :  STD_LOGIC;
                signal sdram_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_s1_arb_counter_enable :  STD_LOGIC;
                signal sdram_s1_arb_share_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sdram_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sdram_s1_arb_share_set_values :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sdram_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal sdram_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sdram_s1_begins_xfer :  STD_LOGIC;
                signal sdram_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sdram_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_s1_end_xfer :  STD_LOGIC;
                signal sdram_s1_firsttransfer :  STD_LOGIC;
                signal sdram_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_s1_in_a_read_cycle :  STD_LOGIC;
                signal sdram_s1_in_a_write_cycle :  STD_LOGIC;
                signal sdram_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal sdram_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sdram_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal sdram_s1_reg_firsttransfer :  STD_LOGIC;
                signal sdram_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sdram_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sdram_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sdram_s1_waits_for_read :  STD_LOGIC;
                signal sdram_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_sdram_s1_from_niosII_system_burst_10_downstream :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal shifted_address_to_sdram_s1_from_niosII_system_burst_11_downstream :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal wait_for_sdram_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sdram_s1_end_xfer;
    end if;

  end process;

  sdram_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_niosII_system_burst_10_downstream_qualified_request_sdram_s1 OR internal_niosII_system_burst_11_downstream_qualified_request_sdram_s1));
  --assign sdram_s1_readdata_from_sa = sdram_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_s1_readdata_from_sa <= sdram_s1_readdata;
  internal_niosII_system_burst_10_downstream_requests_sdram_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_10_downstream_read OR niosII_system_burst_10_downstream_write)))))));
  --assign sdram_s1_waitrequest_from_sa = sdram_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_sdram_s1_waitrequest_from_sa <= sdram_s1_waitrequest;
  --assign sdram_s1_readdatavalid_from_sa = sdram_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_s1_readdatavalid_from_sa <= sdram_s1_readdatavalid;
  --sdram_s1_arb_share_counter set values, which is an e_mux
  sdram_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_10_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_10_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_11_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_11_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_10_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_10_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_11_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_11_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001"))))), 5);
  --sdram_s1_non_bursting_master_requests mux, which is an e_mux
  sdram_s1_non_bursting_master_requests <= std_logic'('0');
  --sdram_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sdram_s1_any_bursting_master_saved_grant <= ((niosII_system_burst_10_downstream_saved_grant_sdram_s1 OR niosII_system_burst_11_downstream_saved_grant_sdram_s1) OR niosII_system_burst_10_downstream_saved_grant_sdram_s1) OR niosII_system_burst_11_downstream_saved_grant_sdram_s1;
  --sdram_s1_arb_share_counter_next_value assignment, which is an e_assign
  sdram_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sdram_s1_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (sdram_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sdram_s1_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (sdram_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 5);
  --sdram_s1_allgrants all slave grants, which is an e_mux
  sdram_s1_allgrants <= (((or_reduce(sdram_s1_grant_vector)) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector));
  --sdram_s1_end_xfer assignment, which is an e_assign
  sdram_s1_end_xfer <= NOT ((sdram_s1_waits_for_read OR sdram_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sdram_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sdram_s1 <= sdram_s1_end_xfer AND (((NOT sdram_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sdram_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sdram_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sdram_s1 AND sdram_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sdram_s1 AND NOT sdram_s1_non_bursting_master_requests));
  --sdram_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_arb_share_counter <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_arb_counter_enable) = '1' then 
        sdram_s1_arb_share_counter <= sdram_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sdram_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(sdram_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_sdram_s1)) OR ((end_xfer_arb_share_counter_term_sdram_s1 AND NOT sdram_s1_non_bursting_master_requests)))) = '1' then 
        sdram_s1_slavearbiterlockenable <= or_reduce(sdram_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_10/downstream sdram/s1 arbiterlock, which is an e_assign
  niosII_system_burst_10_downstream_arbiterlock <= sdram_s1_slavearbiterlockenable AND niosII_system_burst_10_downstream_continuerequest;
  --sdram_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sdram_s1_slavearbiterlockenable2 <= or_reduce(sdram_s1_arb_share_counter_next_value);
  --niosII_system_burst_10/downstream sdram/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_10_downstream_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND niosII_system_burst_10_downstream_continuerequest;
  --niosII_system_burst_11/downstream sdram/s1 arbiterlock, which is an e_assign
  niosII_system_burst_11_downstream_arbiterlock <= sdram_s1_slavearbiterlockenable AND niosII_system_burst_11_downstream_continuerequest;
  --niosII_system_burst_11/downstream sdram/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_11_downstream_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND niosII_system_burst_11_downstream_continuerequest;
  --niosII_system_burst_11/downstream granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_niosII_system_burst_11_downstream_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_niosII_system_burst_11_downstream_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(niosII_system_burst_11_downstream_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_11_downstream_granted_slave_sdram_s1))))));
    end if;

  end process;

  --niosII_system_burst_11_downstream_continuerequest continued request, which is an e_mux
  niosII_system_burst_11_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_11_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --sdram_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  sdram_s1_any_continuerequest <= niosII_system_burst_11_downstream_continuerequest OR niosII_system_burst_10_downstream_continuerequest;
  internal_niosII_system_burst_10_downstream_qualified_request_sdram_s1 <= internal_niosII_system_burst_10_downstream_requests_sdram_s1 AND NOT ((((niosII_system_burst_10_downstream_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_10_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_10_downstream_latency_counter)))))))))) OR niosII_system_burst_11_downstream_arbiterlock));
  --unique name for sdram_s1_move_on_to_next_transaction, which is an e_assign
  sdram_s1_move_on_to_next_transaction <= sdram_s1_readdatavalid_from_sa;
  --rdv_fifo_for_niosII_system_burst_10_downstream_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_niosII_system_burst_10_downstream_to_sdram_s1 : rdv_fifo_for_niosII_system_burst_10_downstream_to_sdram_s1_module
    port map(
      data_out => niosII_system_burst_10_downstream_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => niosII_system_burst_10_downstream_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input132,
      clk => clk,
      data_in => internal_niosII_system_burst_10_downstream_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input133,
      write => module_input134
    );

  module_input132 <= std_logic'('0');
  module_input133 <= std_logic'('0');
  module_input134 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  niosII_system_burst_10_downstream_read_data_valid_sdram_s1_shift_register <= NOT niosII_system_burst_10_downstream_rdv_fifo_empty_sdram_s1;
  --local readdatavalid niosII_system_burst_10_downstream_read_data_valid_sdram_s1, which is an e_mux
  niosII_system_burst_10_downstream_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND niosII_system_burst_10_downstream_rdv_fifo_output_from_sdram_s1)) AND NOT niosII_system_burst_10_downstream_rdv_fifo_empty_sdram_s1;
  --sdram_s1_writedata mux, which is an e_mux
  sdram_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_10_downstream_granted_sdram_s1)) = '1'), niosII_system_burst_10_downstream_writedata, niosII_system_burst_11_downstream_writedata);
  internal_niosII_system_burst_11_downstream_requests_sdram_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_11_downstream_read OR niosII_system_burst_11_downstream_write)))))));
  --niosII_system_burst_10/downstream granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_niosII_system_burst_10_downstream_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_niosII_system_burst_10_downstream_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(niosII_system_burst_10_downstream_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_10_downstream_granted_slave_sdram_s1))))));
    end if;

  end process;

  --niosII_system_burst_10_downstream_continuerequest continued request, which is an e_mux
  niosII_system_burst_10_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_10_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  internal_niosII_system_burst_11_downstream_qualified_request_sdram_s1 <= internal_niosII_system_burst_11_downstream_requests_sdram_s1 AND NOT ((((niosII_system_burst_11_downstream_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_11_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_11_downstream_latency_counter)))))))))) OR niosII_system_burst_10_downstream_arbiterlock));
  --rdv_fifo_for_niosII_system_burst_11_downstream_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_niosII_system_burst_11_downstream_to_sdram_s1 : rdv_fifo_for_niosII_system_burst_11_downstream_to_sdram_s1_module
    port map(
      data_out => niosII_system_burst_11_downstream_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => niosII_system_burst_11_downstream_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input135,
      clk => clk,
      data_in => internal_niosII_system_burst_11_downstream_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input136,
      write => module_input137
    );

  module_input135 <= std_logic'('0');
  module_input136 <= std_logic'('0');
  module_input137 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  niosII_system_burst_11_downstream_read_data_valid_sdram_s1_shift_register <= NOT niosII_system_burst_11_downstream_rdv_fifo_empty_sdram_s1;
  --local readdatavalid niosII_system_burst_11_downstream_read_data_valid_sdram_s1, which is an e_mux
  niosII_system_burst_11_downstream_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND niosII_system_burst_11_downstream_rdv_fifo_output_from_sdram_s1)) AND NOT niosII_system_burst_11_downstream_rdv_fifo_empty_sdram_s1;
  --allow new arb cycle for sdram/s1, which is an e_assign
  sdram_s1_allow_new_arb_cycle <= NOT niosII_system_burst_10_downstream_arbiterlock AND NOT niosII_system_burst_11_downstream_arbiterlock;
  --niosII_system_burst_11/downstream assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(0) <= internal_niosII_system_burst_11_downstream_qualified_request_sdram_s1;
  --niosII_system_burst_11/downstream grant sdram/s1, which is an e_assign
  internal_niosII_system_burst_11_downstream_granted_sdram_s1 <= sdram_s1_grant_vector(0);
  --niosII_system_burst_11/downstream saved-grant sdram/s1, which is an e_assign
  niosII_system_burst_11_downstream_saved_grant_sdram_s1 <= sdram_s1_arb_winner(0);
  --niosII_system_burst_10/downstream assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(1) <= internal_niosII_system_burst_10_downstream_qualified_request_sdram_s1;
  --niosII_system_burst_10/downstream grant sdram/s1, which is an e_assign
  internal_niosII_system_burst_10_downstream_granted_sdram_s1 <= sdram_s1_grant_vector(1);
  --niosII_system_burst_10/downstream saved-grant sdram/s1, which is an e_assign
  niosII_system_burst_10_downstream_saved_grant_sdram_s1 <= sdram_s1_arb_winner(1);
  --sdram/s1 chosen-master double-vector, which is an e_assign
  sdram_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((sdram_s1_master_qreq_vector & sdram_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT sdram_s1_master_qreq_vector & NOT sdram_s1_master_qreq_vector))) + (std_logic_vector'("000") & (sdram_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  sdram_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((sdram_s1_allow_new_arb_cycle AND or_reduce(sdram_s1_grant_vector)))) = '1'), sdram_s1_grant_vector, sdram_s1_saved_chosen_master_vector);
  --saved sdram_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_allow_new_arb_cycle) = '1' then 
        sdram_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(sdram_s1_grant_vector)) = '1'), sdram_s1_grant_vector, sdram_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  sdram_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(1) OR sdram_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(0) OR sdram_s1_chosen_master_double_vector(2)))));
  --sdram/s1 chosen master rotated left, which is an e_assign
  sdram_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(sdram_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(sdram_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --sdram/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(sdram_s1_grant_vector)) = '1' then 
        sdram_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(sdram_s1_end_xfer) = '1'), sdram_s1_chosen_master_rot_left, sdram_s1_grant_vector);
      end if;
    end if;

  end process;

  --sdram_s1_reset_n assignment, which is an e_assign
  sdram_s1_reset_n <= reset_n;
  sdram_s1_chipselect <= internal_niosII_system_burst_10_downstream_granted_sdram_s1 OR internal_niosII_system_burst_11_downstream_granted_sdram_s1;
  --sdram_s1_firsttransfer first transaction, which is an e_assign
  sdram_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sdram_s1_begins_xfer) = '1'), sdram_s1_unreg_firsttransfer, sdram_s1_reg_firsttransfer);
  --sdram_s1_unreg_firsttransfer first transaction, which is an e_assign
  sdram_s1_unreg_firsttransfer <= NOT ((sdram_s1_slavearbiterlockenable AND sdram_s1_any_continuerequest));
  --sdram_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_begins_xfer) = '1' then 
        sdram_s1_reg_firsttransfer <= sdram_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sdram_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sdram_s1_beginbursttransfer_internal <= sdram_s1_begins_xfer;
  --sdram_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  sdram_s1_arbitration_holdoff_internal <= sdram_s1_begins_xfer AND sdram_s1_firsttransfer;
  --~sdram_s1_read_n assignment, which is an e_mux
  sdram_s1_read_n <= NOT ((((internal_niosII_system_burst_10_downstream_granted_sdram_s1 AND niosII_system_burst_10_downstream_read)) OR ((internal_niosII_system_burst_11_downstream_granted_sdram_s1 AND niosII_system_burst_11_downstream_read))));
  --~sdram_s1_write_n assignment, which is an e_mux
  sdram_s1_write_n <= NOT ((((internal_niosII_system_burst_10_downstream_granted_sdram_s1 AND niosII_system_burst_10_downstream_write)) OR ((internal_niosII_system_burst_11_downstream_granted_sdram_s1 AND niosII_system_burst_11_downstream_write))));
  shifted_address_to_sdram_s1_from_niosII_system_burst_10_downstream <= niosII_system_burst_10_downstream_address_to_slave;
  --sdram_s1_address mux, which is an e_mux
  sdram_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_10_downstream_granted_sdram_s1)) = '1'), (A_SRL(shifted_address_to_sdram_s1_from_niosII_system_burst_10_downstream,std_logic_vector'("00000000000000000000000000000001"))), (A_SRL(shifted_address_to_sdram_s1_from_niosII_system_burst_11_downstream,std_logic_vector'("00000000000000000000000000000001")))), 22);
  shifted_address_to_sdram_s1_from_niosII_system_burst_11_downstream <= niosII_system_burst_11_downstream_address_to_slave;
  --d1_sdram_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sdram_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sdram_s1_end_xfer <= sdram_s1_end_xfer;
    end if;

  end process;

  --sdram_s1_waits_for_read in a cycle, which is an e_mux
  sdram_s1_waits_for_read <= sdram_s1_in_a_read_cycle AND internal_sdram_s1_waitrequest_from_sa;
  --sdram_s1_in_a_read_cycle assignment, which is an e_assign
  sdram_s1_in_a_read_cycle <= ((internal_niosII_system_burst_10_downstream_granted_sdram_s1 AND niosII_system_burst_10_downstream_read)) OR ((internal_niosII_system_burst_11_downstream_granted_sdram_s1 AND niosII_system_burst_11_downstream_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sdram_s1_in_a_read_cycle;
  --sdram_s1_waits_for_write in a cycle, which is an e_mux
  sdram_s1_waits_for_write <= sdram_s1_in_a_write_cycle AND internal_sdram_s1_waitrequest_from_sa;
  --sdram_s1_in_a_write_cycle assignment, which is an e_assign
  sdram_s1_in_a_write_cycle <= ((internal_niosII_system_burst_10_downstream_granted_sdram_s1 AND niosII_system_burst_10_downstream_write)) OR ((internal_niosII_system_burst_11_downstream_granted_sdram_s1 AND niosII_system_burst_11_downstream_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sdram_s1_in_a_write_cycle;
  wait_for_sdram_s1_counter <= std_logic'('0');
  --~sdram_s1_byteenable_n byte enable port mux, which is an e_mux
  sdram_s1_byteenable_n <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_10_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_10_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_11_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_11_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))))), 2);
  --vhdl renameroo for output signals
  niosII_system_burst_10_downstream_granted_sdram_s1 <= internal_niosII_system_burst_10_downstream_granted_sdram_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_10_downstream_qualified_request_sdram_s1 <= internal_niosII_system_burst_10_downstream_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_10_downstream_requests_sdram_s1 <= internal_niosII_system_burst_10_downstream_requests_sdram_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_11_downstream_granted_sdram_s1 <= internal_niosII_system_burst_11_downstream_granted_sdram_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_11_downstream_qualified_request_sdram_s1 <= internal_niosII_system_burst_11_downstream_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_11_downstream_requests_sdram_s1 <= internal_niosII_system_burst_11_downstream_requests_sdram_s1;
  --vhdl renameroo for output signals
  sdram_s1_waitrequest_from_sa <= internal_sdram_s1_waitrequest_from_sa;
--synthesis translate_off
    --sdram/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_10/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line192 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_10_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_10_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line192, now);
          write(write_line192, string'(": "));
          write(write_line192, string'("niosII_system_burst_10/downstream drove 0 on its 'arbitrationshare' port while accessing slave sdram/s1"));
          write(output, write_line192.all);
          deallocate (write_line192);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_10/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line193 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_10_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_10_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line193, now);
          write(write_line193, string'(": "));
          write(write_line193, string'("niosII_system_burst_10/downstream drove 0 on its 'burstcount' port while accessing slave sdram/s1"));
          write(output, write_line193.all);
          deallocate (write_line193);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_11/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line194 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_11_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_11_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line194, now);
          write(write_line194, string'(": "));
          write(write_line194, string'("niosII_system_burst_11/downstream drove 0 on its 'arbitrationshare' port while accessing slave sdram/s1"));
          write(output, write_line194.all);
          deallocate (write_line194);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_11/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line195 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_11_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_11_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line195, now);
          write(write_line195, string'(": "));
          write(write_line195, string'("niosII_system_burst_11/downstream drove 0 on its 'burstcount' port while accessing slave sdram/s1"));
          write(output, write_line195.all);
          deallocate (write_line195);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line196 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_10_downstream_granted_sdram_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_11_downstream_granted_sdram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line196, now);
          write(write_line196, string'(": "));
          write(write_line196, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line196.all);
          deallocate (write_line196);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line197 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(niosII_system_burst_10_downstream_saved_grant_sdram_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(niosII_system_burst_11_downstream_saved_grant_sdram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line197, now);
          write(write_line197, string'(": "));
          write(write_line197, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line197.all);
          deallocate (write_line197);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity seven_seg_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_14_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_14_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_14_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_14_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal seven_seg_pio_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal d1_seven_seg_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 : OUT STD_LOGIC;
                 signal seven_seg_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal seven_seg_pio_s1_chipselect : OUT STD_LOGIC;
                 signal seven_seg_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal seven_seg_pio_s1_reset_n : OUT STD_LOGIC;
                 signal seven_seg_pio_s1_write_n : OUT STD_LOGIC;
                 signal seven_seg_pio_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity seven_seg_pio_s1_arbitrator;


architecture europa of seven_seg_pio_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_seven_seg_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_saved_grant_seven_seg_pio_s1 :  STD_LOGIC;
                signal seven_seg_pio_s1_allgrants :  STD_LOGIC;
                signal seven_seg_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal seven_seg_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal seven_seg_pio_s1_any_continuerequest :  STD_LOGIC;
                signal seven_seg_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal seven_seg_pio_s1_arb_share_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal seven_seg_pio_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal seven_seg_pio_s1_arb_share_set_values :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal seven_seg_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal seven_seg_pio_s1_begins_xfer :  STD_LOGIC;
                signal seven_seg_pio_s1_end_xfer :  STD_LOGIC;
                signal seven_seg_pio_s1_firsttransfer :  STD_LOGIC;
                signal seven_seg_pio_s1_grant_vector :  STD_LOGIC;
                signal seven_seg_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal seven_seg_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal seven_seg_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal seven_seg_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal seven_seg_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal seven_seg_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal seven_seg_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal seven_seg_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal seven_seg_pio_s1_waits_for_read :  STD_LOGIC;
                signal seven_seg_pio_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_seven_seg_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT seven_seg_pio_s1_end_xfer;
    end if;

  end process;

  seven_seg_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1);
  --assign seven_seg_pio_s1_readdata_from_sa = seven_seg_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  seven_seg_pio_s1_readdata_from_sa <= seven_seg_pio_s1_readdata;
  internal_niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_14_downstream_read OR niosII_system_burst_14_downstream_write)))))));
  --seven_seg_pio_s1_arb_share_counter set values, which is an e_mux
  seven_seg_pio_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_14_downstream_granted_seven_seg_pio_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_14_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --seven_seg_pio_s1_non_bursting_master_requests mux, which is an e_mux
  seven_seg_pio_s1_non_bursting_master_requests <= std_logic'('0');
  --seven_seg_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  seven_seg_pio_s1_any_bursting_master_saved_grant <= niosII_system_burst_14_downstream_saved_grant_seven_seg_pio_s1;
  --seven_seg_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  seven_seg_pio_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(seven_seg_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (seven_seg_pio_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(seven_seg_pio_s1_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (seven_seg_pio_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 5);
  --seven_seg_pio_s1_allgrants all slave grants, which is an e_mux
  seven_seg_pio_s1_allgrants <= seven_seg_pio_s1_grant_vector;
  --seven_seg_pio_s1_end_xfer assignment, which is an e_assign
  seven_seg_pio_s1_end_xfer <= NOT ((seven_seg_pio_s1_waits_for_read OR seven_seg_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_seven_seg_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_seven_seg_pio_s1 <= seven_seg_pio_s1_end_xfer AND (((NOT seven_seg_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --seven_seg_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  seven_seg_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_seven_seg_pio_s1 AND seven_seg_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_seven_seg_pio_s1 AND NOT seven_seg_pio_s1_non_bursting_master_requests));
  --seven_seg_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      seven_seg_pio_s1_arb_share_counter <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(seven_seg_pio_s1_arb_counter_enable) = '1' then 
        seven_seg_pio_s1_arb_share_counter <= seven_seg_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --seven_seg_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      seven_seg_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((seven_seg_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_seven_seg_pio_s1)) OR ((end_xfer_arb_share_counter_term_seven_seg_pio_s1 AND NOT seven_seg_pio_s1_non_bursting_master_requests)))) = '1' then 
        seven_seg_pio_s1_slavearbiterlockenable <= or_reduce(seven_seg_pio_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_14/downstream seven_seg_pio/s1 arbiterlock, which is an e_assign
  niosII_system_burst_14_downstream_arbiterlock <= seven_seg_pio_s1_slavearbiterlockenable AND niosII_system_burst_14_downstream_continuerequest;
  --seven_seg_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  seven_seg_pio_s1_slavearbiterlockenable2 <= or_reduce(seven_seg_pio_s1_arb_share_counter_next_value);
  --niosII_system_burst_14/downstream seven_seg_pio/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_14_downstream_arbiterlock2 <= seven_seg_pio_s1_slavearbiterlockenable2 AND niosII_system_burst_14_downstream_continuerequest;
  --seven_seg_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  seven_seg_pio_s1_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_14_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_14_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 <= internal_niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 AND NOT ((niosII_system_burst_14_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_14_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1, which is an e_mux
  niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1 <= (internal_niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 AND niosII_system_burst_14_downstream_read) AND NOT seven_seg_pio_s1_waits_for_read;
  --seven_seg_pio_s1_writedata mux, which is an e_mux
  seven_seg_pio_s1_writedata <= niosII_system_burst_14_downstream_writedata;
  --master is always granted when requested
  internal_niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 <= internal_niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1;
  --niosII_system_burst_14/downstream saved-grant seven_seg_pio/s1, which is an e_assign
  niosII_system_burst_14_downstream_saved_grant_seven_seg_pio_s1 <= internal_niosII_system_burst_14_downstream_requests_seven_seg_pio_s1;
  --allow new arb cycle for seven_seg_pio/s1, which is an e_assign
  seven_seg_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  seven_seg_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  seven_seg_pio_s1_master_qreq_vector <= std_logic'('1');
  --seven_seg_pio_s1_reset_n assignment, which is an e_assign
  seven_seg_pio_s1_reset_n <= reset_n;
  seven_seg_pio_s1_chipselect <= internal_niosII_system_burst_14_downstream_granted_seven_seg_pio_s1;
  --seven_seg_pio_s1_firsttransfer first transaction, which is an e_assign
  seven_seg_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(seven_seg_pio_s1_begins_xfer) = '1'), seven_seg_pio_s1_unreg_firsttransfer, seven_seg_pio_s1_reg_firsttransfer);
  --seven_seg_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  seven_seg_pio_s1_unreg_firsttransfer <= NOT ((seven_seg_pio_s1_slavearbiterlockenable AND seven_seg_pio_s1_any_continuerequest));
  --seven_seg_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      seven_seg_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(seven_seg_pio_s1_begins_xfer) = '1' then 
        seven_seg_pio_s1_reg_firsttransfer <= seven_seg_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --seven_seg_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  seven_seg_pio_s1_beginbursttransfer_internal <= seven_seg_pio_s1_begins_xfer;
  --~seven_seg_pio_s1_write_n assignment, which is an e_mux
  seven_seg_pio_s1_write_n <= NOT ((internal_niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 AND niosII_system_burst_14_downstream_write));
  --seven_seg_pio_s1_address mux, which is an e_mux
  seven_seg_pio_s1_address <= niosII_system_burst_14_downstream_nativeaddress (1 DOWNTO 0);
  --d1_seven_seg_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_seven_seg_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_seven_seg_pio_s1_end_xfer <= seven_seg_pio_s1_end_xfer;
    end if;

  end process;

  --seven_seg_pio_s1_waits_for_read in a cycle, which is an e_mux
  seven_seg_pio_s1_waits_for_read <= seven_seg_pio_s1_in_a_read_cycle AND seven_seg_pio_s1_begins_xfer;
  --seven_seg_pio_s1_in_a_read_cycle assignment, which is an e_assign
  seven_seg_pio_s1_in_a_read_cycle <= internal_niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 AND niosII_system_burst_14_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= seven_seg_pio_s1_in_a_read_cycle;
  --seven_seg_pio_s1_waits_for_write in a cycle, which is an e_mux
  seven_seg_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(seven_seg_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --seven_seg_pio_s1_in_a_write_cycle assignment, which is an e_assign
  seven_seg_pio_s1_in_a_write_cycle <= internal_niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 AND niosII_system_burst_14_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= seven_seg_pio_s1_in_a_write_cycle;
  wait_for_seven_seg_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 <= internal_niosII_system_burst_14_downstream_granted_seven_seg_pio_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 <= internal_niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 <= internal_niosII_system_burst_14_downstream_requests_seven_seg_pio_s1;
--synthesis translate_off
    --seven_seg_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_14/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line198 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_14_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line198, now);
          write(write_line198, string'(": "));
          write(write_line198, string'("niosII_system_burst_14/downstream drove 0 on its 'arbitrationshare' port while accessing slave seven_seg_pio/s1"));
          write(output, write_line198.all);
          deallocate (write_line198);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_14/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line199 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_14_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line199, now);
          write(write_line199, string'(": "));
          write(write_line199, string'("niosII_system_burst_14/downstream drove 0 on its 'burstcount' port while accessing slave seven_seg_pio/s1"));
          write(output, write_line199.all);
          deallocate (write_line199);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity switch_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_9_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal niosII_system_burst_9_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_9_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_9_downstream_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal switch_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- outputs:
                 signal d1_switch_s1_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_9_downstream_granted_switch_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_9_downstream_qualified_request_switch_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_9_downstream_read_data_valid_switch_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_9_downstream_requests_switch_s1 : OUT STD_LOGIC;
                 signal switch_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal switch_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal switch_s1_reset_n : OUT STD_LOGIC
              );
end entity switch_s1_arbitrator;


architecture europa of switch_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_switch_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_9_downstream_granted_switch_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_9_downstream_qualified_request_switch_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_9_downstream_requests_switch_s1 :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_saved_grant_switch_s1 :  STD_LOGIC;
                signal switch_s1_allgrants :  STD_LOGIC;
                signal switch_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal switch_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal switch_s1_any_continuerequest :  STD_LOGIC;
                signal switch_s1_arb_counter_enable :  STD_LOGIC;
                signal switch_s1_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal switch_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal switch_s1_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal switch_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal switch_s1_begins_xfer :  STD_LOGIC;
                signal switch_s1_end_xfer :  STD_LOGIC;
                signal switch_s1_firsttransfer :  STD_LOGIC;
                signal switch_s1_grant_vector :  STD_LOGIC;
                signal switch_s1_in_a_read_cycle :  STD_LOGIC;
                signal switch_s1_in_a_write_cycle :  STD_LOGIC;
                signal switch_s1_master_qreq_vector :  STD_LOGIC;
                signal switch_s1_non_bursting_master_requests :  STD_LOGIC;
                signal switch_s1_reg_firsttransfer :  STD_LOGIC;
                signal switch_s1_slavearbiterlockenable :  STD_LOGIC;
                signal switch_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal switch_s1_unreg_firsttransfer :  STD_LOGIC;
                signal switch_s1_waits_for_read :  STD_LOGIC;
                signal switch_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_switch_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT switch_s1_end_xfer;
    end if;

  end process;

  switch_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_9_downstream_qualified_request_switch_s1);
  --assign switch_s1_readdata_from_sa = switch_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  switch_s1_readdata_from_sa <= switch_s1_readdata;
  internal_niosII_system_burst_9_downstream_requests_switch_s1 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_9_downstream_read OR niosII_system_burst_9_downstream_write))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_9_downstream_read)))));
  --switch_s1_arb_share_counter set values, which is an e_mux
  switch_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_9_downstream_granted_switch_s1)) = '1'), (std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_9_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 6);
  --switch_s1_non_bursting_master_requests mux, which is an e_mux
  switch_s1_non_bursting_master_requests <= std_logic'('0');
  --switch_s1_any_bursting_master_saved_grant mux, which is an e_mux
  switch_s1_any_bursting_master_saved_grant <= niosII_system_burst_9_downstream_saved_grant_switch_s1;
  --switch_s1_arb_share_counter_next_value assignment, which is an e_assign
  switch_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(switch_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (switch_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(switch_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (switch_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --switch_s1_allgrants all slave grants, which is an e_mux
  switch_s1_allgrants <= switch_s1_grant_vector;
  --switch_s1_end_xfer assignment, which is an e_assign
  switch_s1_end_xfer <= NOT ((switch_s1_waits_for_read OR switch_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_switch_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_switch_s1 <= switch_s1_end_xfer AND (((NOT switch_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --switch_s1_arb_share_counter arbitration counter enable, which is an e_assign
  switch_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_switch_s1 AND switch_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_switch_s1 AND NOT switch_s1_non_bursting_master_requests));
  --switch_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      switch_s1_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(switch_s1_arb_counter_enable) = '1' then 
        switch_s1_arb_share_counter <= switch_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --switch_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      switch_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((switch_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_switch_s1)) OR ((end_xfer_arb_share_counter_term_switch_s1 AND NOT switch_s1_non_bursting_master_requests)))) = '1' then 
        switch_s1_slavearbiterlockenable <= or_reduce(switch_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_9/downstream switch/s1 arbiterlock, which is an e_assign
  niosII_system_burst_9_downstream_arbiterlock <= switch_s1_slavearbiterlockenable AND niosII_system_burst_9_downstream_continuerequest;
  --switch_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  switch_s1_slavearbiterlockenable2 <= or_reduce(switch_s1_arb_share_counter_next_value);
  --niosII_system_burst_9/downstream switch/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_9_downstream_arbiterlock2 <= switch_s1_slavearbiterlockenable2 AND niosII_system_burst_9_downstream_continuerequest;
  --switch_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  switch_s1_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_9_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_9_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_9_downstream_qualified_request_switch_s1 <= internal_niosII_system_burst_9_downstream_requests_switch_s1 AND NOT ((niosII_system_burst_9_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_9_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_9_downstream_read_data_valid_switch_s1, which is an e_mux
  niosII_system_burst_9_downstream_read_data_valid_switch_s1 <= (internal_niosII_system_burst_9_downstream_granted_switch_s1 AND niosII_system_burst_9_downstream_read) AND NOT switch_s1_waits_for_read;
  --master is always granted when requested
  internal_niosII_system_burst_9_downstream_granted_switch_s1 <= internal_niosII_system_burst_9_downstream_qualified_request_switch_s1;
  --niosII_system_burst_9/downstream saved-grant switch/s1, which is an e_assign
  niosII_system_burst_9_downstream_saved_grant_switch_s1 <= internal_niosII_system_burst_9_downstream_requests_switch_s1;
  --allow new arb cycle for switch/s1, which is an e_assign
  switch_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  switch_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  switch_s1_master_qreq_vector <= std_logic'('1');
  --switch_s1_reset_n assignment, which is an e_assign
  switch_s1_reset_n <= reset_n;
  --switch_s1_firsttransfer first transaction, which is an e_assign
  switch_s1_firsttransfer <= A_WE_StdLogic((std_logic'(switch_s1_begins_xfer) = '1'), switch_s1_unreg_firsttransfer, switch_s1_reg_firsttransfer);
  --switch_s1_unreg_firsttransfer first transaction, which is an e_assign
  switch_s1_unreg_firsttransfer <= NOT ((switch_s1_slavearbiterlockenable AND switch_s1_any_continuerequest));
  --switch_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      switch_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(switch_s1_begins_xfer) = '1' then 
        switch_s1_reg_firsttransfer <= switch_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --switch_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  switch_s1_beginbursttransfer_internal <= switch_s1_begins_xfer;
  --switch_s1_address mux, which is an e_mux
  switch_s1_address <= niosII_system_burst_9_downstream_nativeaddress;
  --d1_switch_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_switch_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_switch_s1_end_xfer <= switch_s1_end_xfer;
    end if;

  end process;

  --switch_s1_waits_for_read in a cycle, which is an e_mux
  switch_s1_waits_for_read <= switch_s1_in_a_read_cycle AND switch_s1_begins_xfer;
  --switch_s1_in_a_read_cycle assignment, which is an e_assign
  switch_s1_in_a_read_cycle <= internal_niosII_system_burst_9_downstream_granted_switch_s1 AND niosII_system_burst_9_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= switch_s1_in_a_read_cycle;
  --switch_s1_waits_for_write in a cycle, which is an e_mux
  switch_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(switch_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --switch_s1_in_a_write_cycle assignment, which is an e_assign
  switch_s1_in_a_write_cycle <= internal_niosII_system_burst_9_downstream_granted_switch_s1 AND niosII_system_burst_9_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= switch_s1_in_a_write_cycle;
  wait_for_switch_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  niosII_system_burst_9_downstream_granted_switch_s1 <= internal_niosII_system_burst_9_downstream_granted_switch_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_9_downstream_qualified_request_switch_s1 <= internal_niosII_system_burst_9_downstream_qualified_request_switch_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_9_downstream_requests_switch_s1 <= internal_niosII_system_burst_9_downstream_requests_switch_s1;
--synthesis translate_off
    --switch/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_9/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line200 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_9_downstream_requests_switch_s1 AND to_std_logic((((std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_9_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line200, now);
          write(write_line200, string'(": "));
          write(write_line200, string'("niosII_system_burst_9/downstream drove 0 on its 'arbitrationshare' port while accessing slave switch/s1"));
          write(output, write_line200.all);
          deallocate (write_line200);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_9/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line201 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_9_downstream_requests_switch_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_9_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line201, now);
          write(write_line201, string'(": "));
          write(write_line201, string'("niosII_system_burst_9/downstream drove 0 on its 'burstcount' port while accessing slave switch/s1"));
          write(output, write_line201.all);
          deallocate (write_line201);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sys_clk_timer_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_5_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_5_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_5_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_timer_s1_irq : IN STD_LOGIC;
                 signal sys_clk_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal d1_sys_clk_timer_s1_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal sys_clk_timer_s1_chipselect : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_irq_from_sa : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sys_clk_timer_s1_reset_n : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_write_n : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sys_clk_timer_s1_arbitrator;


architecture europa of sys_clk_timer_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sys_clk_timer_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_saved_grant_sys_clk_timer_s1 :  STD_LOGIC;
                signal sys_clk_timer_s1_allgrants :  STD_LOGIC;
                signal sys_clk_timer_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sys_clk_timer_s1_any_continuerequest :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_counter_enable :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_share_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sys_clk_timer_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sys_clk_timer_s1_arb_share_set_values :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sys_clk_timer_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sys_clk_timer_s1_begins_xfer :  STD_LOGIC;
                signal sys_clk_timer_s1_end_xfer :  STD_LOGIC;
                signal sys_clk_timer_s1_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_grant_vector :  STD_LOGIC;
                signal sys_clk_timer_s1_in_a_read_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_in_a_write_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_master_qreq_vector :  STD_LOGIC;
                signal sys_clk_timer_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sys_clk_timer_s1_reg_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sys_clk_timer_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sys_clk_timer_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_waits_for_read :  STD_LOGIC;
                signal sys_clk_timer_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_sys_clk_timer_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sys_clk_timer_s1_end_xfer;
    end if;

  end process;

  sys_clk_timer_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1);
  --assign sys_clk_timer_s1_readdata_from_sa = sys_clk_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sys_clk_timer_s1_readdata_from_sa <= sys_clk_timer_s1_readdata;
  internal_niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_5_downstream_read OR niosII_system_burst_5_downstream_write)))))));
  --sys_clk_timer_s1_arb_share_counter set values, which is an e_mux
  sys_clk_timer_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_5_downstream_granted_sys_clk_timer_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_5_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --sys_clk_timer_s1_non_bursting_master_requests mux, which is an e_mux
  sys_clk_timer_s1_non_bursting_master_requests <= std_logic'('0');
  --sys_clk_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sys_clk_timer_s1_any_bursting_master_saved_grant <= niosII_system_burst_5_downstream_saved_grant_sys_clk_timer_s1;
  --sys_clk_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  sys_clk_timer_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sys_clk_timer_s1_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (sys_clk_timer_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sys_clk_timer_s1_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (sys_clk_timer_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 5);
  --sys_clk_timer_s1_allgrants all slave grants, which is an e_mux
  sys_clk_timer_s1_allgrants <= sys_clk_timer_s1_grant_vector;
  --sys_clk_timer_s1_end_xfer assignment, which is an e_assign
  sys_clk_timer_s1_end_xfer <= NOT ((sys_clk_timer_s1_waits_for_read OR sys_clk_timer_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sys_clk_timer_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sys_clk_timer_s1 <= sys_clk_timer_s1_end_xfer AND (((NOT sys_clk_timer_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sys_clk_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sys_clk_timer_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND sys_clk_timer_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND NOT sys_clk_timer_s1_non_bursting_master_requests));
  --sys_clk_timer_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_arb_share_counter <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(sys_clk_timer_s1_arb_counter_enable) = '1' then 
        sys_clk_timer_s1_arb_share_counter <= sys_clk_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sys_clk_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sys_clk_timer_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_sys_clk_timer_s1)) OR ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND NOT sys_clk_timer_s1_non_bursting_master_requests)))) = '1' then 
        sys_clk_timer_s1_slavearbiterlockenable <= or_reduce(sys_clk_timer_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_5/downstream sys_clk_timer/s1 arbiterlock, which is an e_assign
  niosII_system_burst_5_downstream_arbiterlock <= sys_clk_timer_s1_slavearbiterlockenable AND niosII_system_burst_5_downstream_continuerequest;
  --sys_clk_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sys_clk_timer_s1_slavearbiterlockenable2 <= or_reduce(sys_clk_timer_s1_arb_share_counter_next_value);
  --niosII_system_burst_5/downstream sys_clk_timer/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_5_downstream_arbiterlock2 <= sys_clk_timer_s1_slavearbiterlockenable2 AND niosII_system_burst_5_downstream_continuerequest;
  --sys_clk_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  sys_clk_timer_s1_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_5_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_5_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 <= internal_niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 AND NOT ((niosII_system_burst_5_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_5_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1, which is an e_mux
  niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1 <= (internal_niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 AND niosII_system_burst_5_downstream_read) AND NOT sys_clk_timer_s1_waits_for_read;
  --sys_clk_timer_s1_writedata mux, which is an e_mux
  sys_clk_timer_s1_writedata <= niosII_system_burst_5_downstream_writedata;
  --master is always granted when requested
  internal_niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 <= internal_niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1;
  --niosII_system_burst_5/downstream saved-grant sys_clk_timer/s1, which is an e_assign
  niosII_system_burst_5_downstream_saved_grant_sys_clk_timer_s1 <= internal_niosII_system_burst_5_downstream_requests_sys_clk_timer_s1;
  --allow new arb cycle for sys_clk_timer/s1, which is an e_assign
  sys_clk_timer_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sys_clk_timer_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sys_clk_timer_s1_master_qreq_vector <= std_logic'('1');
  --sys_clk_timer_s1_reset_n assignment, which is an e_assign
  sys_clk_timer_s1_reset_n <= reset_n;
  sys_clk_timer_s1_chipselect <= internal_niosII_system_burst_5_downstream_granted_sys_clk_timer_s1;
  --sys_clk_timer_s1_firsttransfer first transaction, which is an e_assign
  sys_clk_timer_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sys_clk_timer_s1_begins_xfer) = '1'), sys_clk_timer_s1_unreg_firsttransfer, sys_clk_timer_s1_reg_firsttransfer);
  --sys_clk_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  sys_clk_timer_s1_unreg_firsttransfer <= NOT ((sys_clk_timer_s1_slavearbiterlockenable AND sys_clk_timer_s1_any_continuerequest));
  --sys_clk_timer_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sys_clk_timer_s1_begins_xfer) = '1' then 
        sys_clk_timer_s1_reg_firsttransfer <= sys_clk_timer_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sys_clk_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sys_clk_timer_s1_beginbursttransfer_internal <= sys_clk_timer_s1_begins_xfer;
  --~sys_clk_timer_s1_write_n assignment, which is an e_mux
  sys_clk_timer_s1_write_n <= NOT ((internal_niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 AND niosII_system_burst_5_downstream_write));
  --sys_clk_timer_s1_address mux, which is an e_mux
  sys_clk_timer_s1_address <= niosII_system_burst_5_downstream_nativeaddress (2 DOWNTO 0);
  --d1_sys_clk_timer_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sys_clk_timer_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sys_clk_timer_s1_end_xfer <= sys_clk_timer_s1_end_xfer;
    end if;

  end process;

  --sys_clk_timer_s1_waits_for_read in a cycle, which is an e_mux
  sys_clk_timer_s1_waits_for_read <= sys_clk_timer_s1_in_a_read_cycle AND sys_clk_timer_s1_begins_xfer;
  --sys_clk_timer_s1_in_a_read_cycle assignment, which is an e_assign
  sys_clk_timer_s1_in_a_read_cycle <= internal_niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 AND niosII_system_burst_5_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sys_clk_timer_s1_in_a_read_cycle;
  --sys_clk_timer_s1_waits_for_write in a cycle, which is an e_mux
  sys_clk_timer_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_timer_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sys_clk_timer_s1_in_a_write_cycle assignment, which is an e_assign
  sys_clk_timer_s1_in_a_write_cycle <= internal_niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 AND niosII_system_burst_5_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sys_clk_timer_s1_in_a_write_cycle;
  wait_for_sys_clk_timer_s1_counter <= std_logic'('0');
  --assign sys_clk_timer_s1_irq_from_sa = sys_clk_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sys_clk_timer_s1_irq_from_sa <= sys_clk_timer_s1_irq;
  --vhdl renameroo for output signals
  niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 <= internal_niosII_system_burst_5_downstream_granted_sys_clk_timer_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 <= internal_niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 <= internal_niosII_system_burst_5_downstream_requests_sys_clk_timer_s1;
--synthesis translate_off
    --sys_clk_timer/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_5/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line202 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_5_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line202, now);
          write(write_line202, string'(": "));
          write(write_line202, string'("niosII_system_burst_5/downstream drove 0 on its 'arbitrationshare' port while accessing slave sys_clk_timer/s1"));
          write(output, write_line202.all);
          deallocate (write_line202);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_5/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line203 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_5_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line203, now);
          write(write_line203, string'(": "));
          write(write_line203, string'("niosII_system_burst_5/downstream drove 0 on its 'burstcount' port while accessing slave sys_clk_timer/s1"));
          write(output, write_line203.all);
          deallocate (write_line203);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sysid_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_4_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_4_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_system_burst_4_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_4_downstream_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_4_downstream_granted_sysid_control_slave : OUT STD_LOGIC;
                 signal niosII_system_burst_4_downstream_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                 signal niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                 signal niosII_system_burst_4_downstream_requests_sysid_control_slave : OUT STD_LOGIC;
                 signal sysid_control_slave_address : OUT STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sysid_control_slave_reset_n : OUT STD_LOGIC
              );
end entity sysid_control_slave_arbitrator;


architecture europa of sysid_control_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sysid_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_4_downstream_granted_sysid_control_slave :  STD_LOGIC;
                signal internal_niosII_system_burst_4_downstream_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal internal_niosII_system_burst_4_downstream_requests_sysid_control_slave :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_saved_grant_sysid_control_slave :  STD_LOGIC;
                signal sysid_control_slave_allgrants :  STD_LOGIC;
                signal sysid_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal sysid_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sysid_control_slave_any_continuerequest :  STD_LOGIC;
                signal sysid_control_slave_arb_counter_enable :  STD_LOGIC;
                signal sysid_control_slave_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sysid_control_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sysid_control_slave_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sysid_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal sysid_control_slave_begins_xfer :  STD_LOGIC;
                signal sysid_control_slave_end_xfer :  STD_LOGIC;
                signal sysid_control_slave_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_grant_vector :  STD_LOGIC;
                signal sysid_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal sysid_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal sysid_control_slave_master_qreq_vector :  STD_LOGIC;
                signal sysid_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal sysid_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal sysid_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_waits_for_read :  STD_LOGIC;
                signal sysid_control_slave_waits_for_write :  STD_LOGIC;
                signal wait_for_sysid_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sysid_control_slave_end_xfer;
    end if;

  end process;

  sysid_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_4_downstream_qualified_request_sysid_control_slave);
  --assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sysid_control_slave_readdata_from_sa <= sysid_control_slave_readdata;
  internal_niosII_system_burst_4_downstream_requests_sysid_control_slave <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_4_downstream_read OR niosII_system_burst_4_downstream_write))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_4_downstream_read)))));
  --sysid_control_slave_arb_share_counter set values, which is an e_mux
  sysid_control_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_4_downstream_granted_sysid_control_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_4_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  sysid_control_slave_non_bursting_master_requests <= std_logic'('0');
  --sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  sysid_control_slave_any_bursting_master_saved_grant <= niosII_system_burst_4_downstream_saved_grant_sysid_control_slave;
  --sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  sysid_control_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sysid_control_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (sysid_control_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sysid_control_slave_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (sysid_control_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --sysid_control_slave_allgrants all slave grants, which is an e_mux
  sysid_control_slave_allgrants <= sysid_control_slave_grant_vector;
  --sysid_control_slave_end_xfer assignment, which is an e_assign
  sysid_control_slave_end_xfer <= NOT ((sysid_control_slave_waits_for_read OR sysid_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sysid_control_slave <= sysid_control_slave_end_xfer AND (((NOT sysid_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  sysid_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sysid_control_slave AND sysid_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests));
  --sysid_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_arb_counter_enable) = '1' then 
        sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sysid_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_sysid_control_slave)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests)))) = '1' then 
        sysid_control_slave_slavearbiterlockenable <= or_reduce(sysid_control_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_4/downstream sysid/control_slave arbiterlock, which is an e_assign
  niosII_system_burst_4_downstream_arbiterlock <= sysid_control_slave_slavearbiterlockenable AND niosII_system_burst_4_downstream_continuerequest;
  --sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sysid_control_slave_slavearbiterlockenable2 <= or_reduce(sysid_control_slave_arb_share_counter_next_value);
  --niosII_system_burst_4/downstream sysid/control_slave arbiterlock2, which is an e_assign
  niosII_system_burst_4_downstream_arbiterlock2 <= sysid_control_slave_slavearbiterlockenable2 AND niosII_system_burst_4_downstream_continuerequest;
  --sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  sysid_control_slave_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_4_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_4_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_4_downstream_qualified_request_sysid_control_slave <= internal_niosII_system_burst_4_downstream_requests_sysid_control_slave AND NOT ((niosII_system_burst_4_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_4_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave, which is an e_mux
  niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave <= (internal_niosII_system_burst_4_downstream_granted_sysid_control_slave AND niosII_system_burst_4_downstream_read) AND NOT sysid_control_slave_waits_for_read;
  --master is always granted when requested
  internal_niosII_system_burst_4_downstream_granted_sysid_control_slave <= internal_niosII_system_burst_4_downstream_qualified_request_sysid_control_slave;
  --niosII_system_burst_4/downstream saved-grant sysid/control_slave, which is an e_assign
  niosII_system_burst_4_downstream_saved_grant_sysid_control_slave <= internal_niosII_system_burst_4_downstream_requests_sysid_control_slave;
  --allow new arb cycle for sysid/control_slave, which is an e_assign
  sysid_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sysid_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sysid_control_slave_master_qreq_vector <= std_logic'('1');
  --sysid_control_slave_reset_n assignment, which is an e_assign
  sysid_control_slave_reset_n <= reset_n;
  --sysid_control_slave_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(sysid_control_slave_begins_xfer) = '1'), sysid_control_slave_unreg_firsttransfer, sysid_control_slave_reg_firsttransfer);
  --sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_unreg_firsttransfer <= NOT ((sysid_control_slave_slavearbiterlockenable AND sysid_control_slave_any_continuerequest));
  --sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_begins_xfer) = '1' then 
        sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sysid_control_slave_beginbursttransfer_internal <= sysid_control_slave_begins_xfer;
  --sysid_control_slave_address mux, which is an e_mux
  sysid_control_slave_address <= niosII_system_burst_4_downstream_nativeaddress(0);
  --d1_sysid_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sysid_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end if;

  end process;

  --sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  sysid_control_slave_waits_for_read <= sysid_control_slave_in_a_read_cycle AND sysid_control_slave_begins_xfer;
  --sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_read_cycle <= internal_niosII_system_burst_4_downstream_granted_sysid_control_slave AND niosII_system_burst_4_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sysid_control_slave_in_a_read_cycle;
  --sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  sysid_control_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_write_cycle <= internal_niosII_system_burst_4_downstream_granted_sysid_control_slave AND niosII_system_burst_4_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sysid_control_slave_in_a_write_cycle;
  wait_for_sysid_control_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  niosII_system_burst_4_downstream_granted_sysid_control_slave <= internal_niosII_system_burst_4_downstream_granted_sysid_control_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_4_downstream_qualified_request_sysid_control_slave <= internal_niosII_system_burst_4_downstream_qualified_request_sysid_control_slave;
  --vhdl renameroo for output signals
  niosII_system_burst_4_downstream_requests_sysid_control_slave <= internal_niosII_system_burst_4_downstream_requests_sysid_control_slave;
--synthesis translate_off
    --sysid/control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_4/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line204 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_4_downstream_requests_sysid_control_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (niosII_system_burst_4_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line204, now);
          write(write_line204, string'(": "));
          write(write_line204, string'("niosII_system_burst_4/downstream drove 0 on its 'arbitrationshare' port while accessing slave sysid/control_slave"));
          write(output, write_line204.all);
          deallocate (write_line204);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_4/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line205 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_4_downstream_requests_sysid_control_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_4_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line205, now);
          write(write_line205, string'(": "));
          write(write_line205, string'("niosII_system_burst_4/downstream drove 0 on its 'burstcount' port while accessing slave sysid/control_slave"));
          write(output, write_line205.all);
          deallocate (write_line205);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity tri_state_bridge_avalon_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_address_to_slave : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal niosII_system_burst_12_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal niosII_system_burst_12_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_byteenable : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_12_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_12_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_13_downstream_address_to_slave : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal niosII_system_burst_13_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal niosII_system_burst_13_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_byteenable : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_13_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_13_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal address_to_the_ext_flash : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal d1_tri_state_bridge_avalon_slave_end_xfer : OUT STD_LOGIC;
                 signal data_to_and_from_the_ext_flash : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal ext_flash_s1_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_system_burst_12_downstream_granted_ext_flash_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_12_downstream_requests_ext_flash_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_13_downstream_granted_ext_flash_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_13_downstream_requests_ext_flash_s1 : OUT STD_LOGIC;
                 signal read_n_to_the_ext_flash : OUT STD_LOGIC;
                 signal select_n_to_the_ext_flash : OUT STD_LOGIC;
                 signal write_n_to_the_ext_flash : OUT STD_LOGIC
              );
end entity tri_state_bridge_avalon_slave_arbitrator;


architecture europa of tri_state_bridge_avalon_slave_arbitrator is
                signal d1_in_a_write_cycle :  STD_LOGIC;
                signal d1_outgoing_data_to_and_from_the_ext_flash :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_tri_state_bridge_avalon_slave :  STD_LOGIC;
                signal ext_flash_s1_counter_load_value :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal ext_flash_s1_in_a_read_cycle :  STD_LOGIC;
                signal ext_flash_s1_in_a_write_cycle :  STD_LOGIC;
                signal ext_flash_s1_pretend_byte_enable :  STD_LOGIC;
                signal ext_flash_s1_wait_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal ext_flash_s1_waits_for_read :  STD_LOGIC;
                signal ext_flash_s1_waits_for_write :  STD_LOGIC;
                signal ext_flash_s1_with_write_latency :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal incoming_data_to_and_from_the_ext_flash :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal incoming_data_to_and_from_the_ext_flash_bit_0_is_x :  STD_LOGIC;
                signal incoming_data_to_and_from_the_ext_flash_bit_1_is_x :  STD_LOGIC;
                signal incoming_data_to_and_from_the_ext_flash_bit_2_is_x :  STD_LOGIC;
                signal incoming_data_to_and_from_the_ext_flash_bit_3_is_x :  STD_LOGIC;
                signal incoming_data_to_and_from_the_ext_flash_bit_4_is_x :  STD_LOGIC;
                signal incoming_data_to_and_from_the_ext_flash_bit_5_is_x :  STD_LOGIC;
                signal incoming_data_to_and_from_the_ext_flash_bit_6_is_x :  STD_LOGIC;
                signal incoming_data_to_and_from_the_ext_flash_bit_7_is_x :  STD_LOGIC;
                signal internal_ext_flash_s1_wait_counter_eq_0 :  STD_LOGIC;
                signal internal_niosII_system_burst_12_downstream_granted_ext_flash_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_12_downstream_requests_ext_flash_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_13_downstream_granted_ext_flash_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_13_downstream_requests_ext_flash_s1 :  STD_LOGIC;
                signal last_cycle_niosII_system_burst_12_downstream_granted_slave_ext_flash_s1 :  STD_LOGIC;
                signal last_cycle_niosII_system_burst_13_downstream_granted_slave_ext_flash_s1 :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register_in :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_saved_grant_ext_flash_s1 :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register_in :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_saved_grant_ext_flash_s1 :  STD_LOGIC;
                signal outgoing_data_to_and_from_the_ext_flash :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_address_to_the_ext_flash :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal p1_niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_read_n_to_the_ext_flash :  STD_LOGIC;
                signal p1_select_n_to_the_ext_flash :  STD_LOGIC;
                signal p1_write_n_to_the_ext_flash :  STD_LOGIC;
                signal time_to_write :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_allgrants :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_any_continuerequest :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tri_state_bridge_avalon_slave_arb_counter_enable :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal tri_state_bridge_avalon_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal tri_state_bridge_avalon_slave_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal tri_state_bridge_avalon_slave_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tri_state_bridge_avalon_slave_arbitration_holdoff_internal :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_begins_xfer :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tri_state_bridge_avalon_slave_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tri_state_bridge_avalon_slave_end_xfer :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_firsttransfer :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tri_state_bridge_avalon_slave_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tri_state_bridge_avalon_slave_non_bursting_master_requests :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_read_pending :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_reg_firsttransfer :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tri_state_bridge_avalon_slave_slavearbiterlockenable :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_unreg_firsttransfer :  STD_LOGIC;
                signal tri_state_bridge_avalon_slave_write_pending :  STD_LOGIC;
                signal wait_for_ext_flash_s1_counter :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of address_to_the_ext_flash : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of d1_in_a_write_cycle : signal is "FAST_OUTPUT_ENABLE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of d1_outgoing_data_to_and_from_the_ext_flash : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of incoming_data_to_and_from_the_ext_flash : signal is "FAST_INPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of read_n_to_the_ext_flash : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of select_n_to_the_ext_flash : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of write_n_to_the_ext_flash : signal is "FAST_OUTPUT_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT tri_state_bridge_avalon_slave_end_xfer;
    end if;

  end process;

  tri_state_bridge_avalon_slave_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 OR internal_niosII_system_burst_13_downstream_qualified_request_ext_flash_s1));
  internal_niosII_system_burst_12_downstream_requests_ext_flash_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_12_downstream_read OR niosII_system_burst_12_downstream_write)))))));
  --~select_n_to_the_ext_flash of type chipselect to ~p1_select_n_to_the_ext_flash, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      select_n_to_the_ext_flash <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      select_n_to_the_ext_flash <= p1_select_n_to_the_ext_flash;
    end if;

  end process;

  tri_state_bridge_avalon_slave_write_pending <= std_logic'('0');
  --tri_state_bridge/avalon_slave read pending calc, which is an e_assign
  tri_state_bridge_avalon_slave_read_pending <= std_logic'('0');
  --tri_state_bridge_avalon_slave_arb_share_counter set values, which is an e_mux
  tri_state_bridge_avalon_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_12_downstream_granted_ext_flash_s1)) = '1'), (std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_12_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_13_downstream_granted_ext_flash_s1)) = '1'), (std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_13_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_12_downstream_granted_ext_flash_s1)) = '1'), (std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_12_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_13_downstream_granted_ext_flash_s1)) = '1'), (std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_13_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001"))))), 6);
  --tri_state_bridge_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  tri_state_bridge_avalon_slave_non_bursting_master_requests <= std_logic'('0');
  --tri_state_bridge_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  tri_state_bridge_avalon_slave_any_bursting_master_saved_grant <= ((niosII_system_burst_12_downstream_saved_grant_ext_flash_s1 OR niosII_system_burst_13_downstream_saved_grant_ext_flash_s1) OR niosII_system_burst_12_downstream_saved_grant_ext_flash_s1) OR niosII_system_burst_13_downstream_saved_grant_ext_flash_s1;
  --tri_state_bridge_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  tri_state_bridge_avalon_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(tri_state_bridge_avalon_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (tri_state_bridge_avalon_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(tri_state_bridge_avalon_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (tri_state_bridge_avalon_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --tri_state_bridge_avalon_slave_allgrants all slave grants, which is an e_mux
  tri_state_bridge_avalon_slave_allgrants <= (((or_reduce(tri_state_bridge_avalon_slave_grant_vector)) OR (or_reduce(tri_state_bridge_avalon_slave_grant_vector))) OR (or_reduce(tri_state_bridge_avalon_slave_grant_vector))) OR (or_reduce(tri_state_bridge_avalon_slave_grant_vector));
  --tri_state_bridge_avalon_slave_end_xfer assignment, which is an e_assign
  tri_state_bridge_avalon_slave_end_xfer <= NOT ((ext_flash_s1_waits_for_read OR ext_flash_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_tri_state_bridge_avalon_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_tri_state_bridge_avalon_slave <= tri_state_bridge_avalon_slave_end_xfer AND (((NOT tri_state_bridge_avalon_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --tri_state_bridge_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  tri_state_bridge_avalon_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_tri_state_bridge_avalon_slave AND tri_state_bridge_avalon_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_tri_state_bridge_avalon_slave AND NOT tri_state_bridge_avalon_slave_non_bursting_master_requests));
  --tri_state_bridge_avalon_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_avalon_slave_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(tri_state_bridge_avalon_slave_arb_counter_enable) = '1' then 
        tri_state_bridge_avalon_slave_arb_share_counter <= tri_state_bridge_avalon_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --tri_state_bridge_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_avalon_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(tri_state_bridge_avalon_slave_master_qreq_vector) AND end_xfer_arb_share_counter_term_tri_state_bridge_avalon_slave)) OR ((end_xfer_arb_share_counter_term_tri_state_bridge_avalon_slave AND NOT tri_state_bridge_avalon_slave_non_bursting_master_requests)))) = '1' then 
        tri_state_bridge_avalon_slave_slavearbiterlockenable <= or_reduce(tri_state_bridge_avalon_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_12/downstream tri_state_bridge/avalon_slave arbiterlock, which is an e_assign
  niosII_system_burst_12_downstream_arbiterlock <= tri_state_bridge_avalon_slave_slavearbiterlockenable AND niosII_system_burst_12_downstream_continuerequest;
  --tri_state_bridge_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  tri_state_bridge_avalon_slave_slavearbiterlockenable2 <= or_reduce(tri_state_bridge_avalon_slave_arb_share_counter_next_value);
  --niosII_system_burst_12/downstream tri_state_bridge/avalon_slave arbiterlock2, which is an e_assign
  niosII_system_burst_12_downstream_arbiterlock2 <= tri_state_bridge_avalon_slave_slavearbiterlockenable2 AND niosII_system_burst_12_downstream_continuerequest;
  --niosII_system_burst_13/downstream tri_state_bridge/avalon_slave arbiterlock, which is an e_assign
  niosII_system_burst_13_downstream_arbiterlock <= tri_state_bridge_avalon_slave_slavearbiterlockenable AND niosII_system_burst_13_downstream_continuerequest;
  --niosII_system_burst_13/downstream tri_state_bridge/avalon_slave arbiterlock2, which is an e_assign
  niosII_system_burst_13_downstream_arbiterlock2 <= tri_state_bridge_avalon_slave_slavearbiterlockenable2 AND niosII_system_burst_13_downstream_continuerequest;
  --niosII_system_burst_13/downstream granted ext_flash/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_niosII_system_burst_13_downstream_granted_slave_ext_flash_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_niosII_system_burst_13_downstream_granted_slave_ext_flash_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(niosII_system_burst_13_downstream_saved_grant_ext_flash_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tri_state_bridge_avalon_slave_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_13_downstream_granted_slave_ext_flash_s1))))));
    end if;

  end process;

  --niosII_system_burst_13_downstream_continuerequest continued request, which is an e_mux
  niosII_system_burst_13_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_13_downstream_granted_slave_ext_flash_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --tri_state_bridge_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  tri_state_bridge_avalon_slave_any_continuerequest <= niosII_system_burst_13_downstream_continuerequest OR niosII_system_burst_12_downstream_continuerequest;
  internal_niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 <= internal_niosII_system_burst_12_downstream_requests_ext_flash_s1 AND NOT (((((niosII_system_burst_12_downstream_read AND ((tri_state_bridge_avalon_slave_write_pending OR (tri_state_bridge_avalon_slave_read_pending))))) OR (((tri_state_bridge_avalon_slave_read_pending) AND niosII_system_burst_12_downstream_write))) OR niosII_system_burst_13_downstream_arbiterlock));
  --niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register_in <= (internal_niosII_system_burst_12_downstream_granted_ext_flash_s1 AND niosII_system_burst_12_downstream_read) AND NOT ext_flash_s1_waits_for_read;
  --shift register p1 niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register <= A_EXT ((niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register & A_ToStdLogicVector(niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register_in)), 2);
  --niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register <= p1_niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register;
    end if;

  end process;

  --local readdatavalid niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1, which is an e_mux
  niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1 <= niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1_shift_register(1);
  --data_to_and_from_the_ext_flash register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      incoming_data_to_and_from_the_ext_flash <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      incoming_data_to_and_from_the_ext_flash <= data_to_and_from_the_ext_flash;
    end if;

  end process;

  --ext_flash_s1_with_write_latency assignment, which is an e_assign
  ext_flash_s1_with_write_latency <= in_a_write_cycle AND ((internal_niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 OR internal_niosII_system_burst_13_downstream_qualified_request_ext_flash_s1));
  --time to write the data, which is an e_mux
  time_to_write <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((ext_flash_s1_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((ext_flash_s1_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), std_logic_vector'("00000000000000000000000000000000"))));
  --d1_outgoing_data_to_and_from_the_ext_flash register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_outgoing_data_to_and_from_the_ext_flash <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      d1_outgoing_data_to_and_from_the_ext_flash <= outgoing_data_to_and_from_the_ext_flash;
    end if;

  end process;

  --write cycle delayed by 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_in_a_write_cycle <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_in_a_write_cycle <= time_to_write;
    end if;

  end process;

  --d1_outgoing_data_to_and_from_the_ext_flash tristate driver, which is an e_assign
  data_to_and_from_the_ext_flash <= A_WE_StdLogicVector((std_logic'((d1_in_a_write_cycle)) = '1'), d1_outgoing_data_to_and_from_the_ext_flash, A_REP(std_logic'('Z'), 8));
  --outgoing_data_to_and_from_the_ext_flash mux, which is an e_mux
  outgoing_data_to_and_from_the_ext_flash <= A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_12_downstream_granted_ext_flash_s1)) = '1'), niosII_system_burst_12_downstream_writedata, niosII_system_burst_13_downstream_writedata);
  internal_niosII_system_burst_13_downstream_requests_ext_flash_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_13_downstream_read OR niosII_system_burst_13_downstream_write)))))));
  --niosII_system_burst_12/downstream granted ext_flash/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_niosII_system_burst_12_downstream_granted_slave_ext_flash_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_niosII_system_burst_12_downstream_granted_slave_ext_flash_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(niosII_system_burst_12_downstream_saved_grant_ext_flash_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tri_state_bridge_avalon_slave_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_12_downstream_granted_slave_ext_flash_s1))))));
    end if;

  end process;

  --niosII_system_burst_12_downstream_continuerequest continued request, which is an e_mux
  niosII_system_burst_12_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_12_downstream_granted_slave_ext_flash_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  internal_niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 <= internal_niosII_system_burst_13_downstream_requests_ext_flash_s1 AND NOT (((((niosII_system_burst_13_downstream_read AND ((tri_state_bridge_avalon_slave_write_pending OR (tri_state_bridge_avalon_slave_read_pending))))) OR (((tri_state_bridge_avalon_slave_read_pending) AND niosII_system_burst_13_downstream_write))) OR niosII_system_burst_12_downstream_arbiterlock));
  --niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register_in <= (internal_niosII_system_burst_13_downstream_granted_ext_flash_s1 AND niosII_system_burst_13_downstream_read) AND NOT ext_flash_s1_waits_for_read;
  --shift register p1 niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register <= A_EXT ((niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register & A_ToStdLogicVector(niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register_in)), 2);
  --niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register <= p1_niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register;
    end if;

  end process;

  --local readdatavalid niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1, which is an e_mux
  niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1 <= niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1_shift_register(1);
  --allow new arb cycle for tri_state_bridge/avalon_slave, which is an e_assign
  tri_state_bridge_avalon_slave_allow_new_arb_cycle <= NOT niosII_system_burst_12_downstream_arbiterlock AND NOT niosII_system_burst_13_downstream_arbiterlock;
  --niosII_system_burst_13/downstream assignment into master qualified-requests vector for ext_flash/s1, which is an e_assign
  tri_state_bridge_avalon_slave_master_qreq_vector(0) <= internal_niosII_system_burst_13_downstream_qualified_request_ext_flash_s1;
  --niosII_system_burst_13/downstream grant ext_flash/s1, which is an e_assign
  internal_niosII_system_burst_13_downstream_granted_ext_flash_s1 <= tri_state_bridge_avalon_slave_grant_vector(0);
  --niosII_system_burst_13/downstream saved-grant ext_flash/s1, which is an e_assign
  niosII_system_burst_13_downstream_saved_grant_ext_flash_s1 <= tri_state_bridge_avalon_slave_arb_winner(0);
  --niosII_system_burst_12/downstream assignment into master qualified-requests vector for ext_flash/s1, which is an e_assign
  tri_state_bridge_avalon_slave_master_qreq_vector(1) <= internal_niosII_system_burst_12_downstream_qualified_request_ext_flash_s1;
  --niosII_system_burst_12/downstream grant ext_flash/s1, which is an e_assign
  internal_niosII_system_burst_12_downstream_granted_ext_flash_s1 <= tri_state_bridge_avalon_slave_grant_vector(1);
  --niosII_system_burst_12/downstream saved-grant ext_flash/s1, which is an e_assign
  niosII_system_burst_12_downstream_saved_grant_ext_flash_s1 <= tri_state_bridge_avalon_slave_arb_winner(1);
  --tri_state_bridge/avalon_slave chosen-master double-vector, which is an e_assign
  tri_state_bridge_avalon_slave_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((tri_state_bridge_avalon_slave_master_qreq_vector & tri_state_bridge_avalon_slave_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT tri_state_bridge_avalon_slave_master_qreq_vector & NOT tri_state_bridge_avalon_slave_master_qreq_vector))) + (std_logic_vector'("000") & (tri_state_bridge_avalon_slave_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  tri_state_bridge_avalon_slave_arb_winner <= A_WE_StdLogicVector((std_logic'(((tri_state_bridge_avalon_slave_allow_new_arb_cycle AND or_reduce(tri_state_bridge_avalon_slave_grant_vector)))) = '1'), tri_state_bridge_avalon_slave_grant_vector, tri_state_bridge_avalon_slave_saved_chosen_master_vector);
  --saved tri_state_bridge_avalon_slave_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_avalon_slave_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(tri_state_bridge_avalon_slave_allow_new_arb_cycle) = '1' then 
        tri_state_bridge_avalon_slave_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(tri_state_bridge_avalon_slave_grant_vector)) = '1'), tri_state_bridge_avalon_slave_grant_vector, tri_state_bridge_avalon_slave_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  tri_state_bridge_avalon_slave_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((tri_state_bridge_avalon_slave_chosen_master_double_vector(1) OR tri_state_bridge_avalon_slave_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((tri_state_bridge_avalon_slave_chosen_master_double_vector(0) OR tri_state_bridge_avalon_slave_chosen_master_double_vector(2)))));
  --tri_state_bridge/avalon_slave chosen master rotated left, which is an e_assign
  tri_state_bridge_avalon_slave_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(tri_state_bridge_avalon_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(tri_state_bridge_avalon_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --tri_state_bridge/avalon_slave's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_avalon_slave_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(tri_state_bridge_avalon_slave_grant_vector)) = '1' then 
        tri_state_bridge_avalon_slave_arb_addend <= A_WE_StdLogicVector((std_logic'(tri_state_bridge_avalon_slave_end_xfer) = '1'), tri_state_bridge_avalon_slave_chosen_master_rot_left, tri_state_bridge_avalon_slave_grant_vector);
      end if;
    end if;

  end process;

  p1_select_n_to_the_ext_flash <= NOT ((internal_niosII_system_burst_12_downstream_granted_ext_flash_s1 OR internal_niosII_system_burst_13_downstream_granted_ext_flash_s1));
  --tri_state_bridge_avalon_slave_firsttransfer first transaction, which is an e_assign
  tri_state_bridge_avalon_slave_firsttransfer <= A_WE_StdLogic((std_logic'(tri_state_bridge_avalon_slave_begins_xfer) = '1'), tri_state_bridge_avalon_slave_unreg_firsttransfer, tri_state_bridge_avalon_slave_reg_firsttransfer);
  --tri_state_bridge_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  tri_state_bridge_avalon_slave_unreg_firsttransfer <= NOT ((tri_state_bridge_avalon_slave_slavearbiterlockenable AND tri_state_bridge_avalon_slave_any_continuerequest));
  --tri_state_bridge_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_avalon_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(tri_state_bridge_avalon_slave_begins_xfer) = '1' then 
        tri_state_bridge_avalon_slave_reg_firsttransfer <= tri_state_bridge_avalon_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --tri_state_bridge_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  tri_state_bridge_avalon_slave_beginbursttransfer_internal <= tri_state_bridge_avalon_slave_begins_xfer;
  --tri_state_bridge_avalon_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  tri_state_bridge_avalon_slave_arbitration_holdoff_internal <= tri_state_bridge_avalon_slave_begins_xfer AND tri_state_bridge_avalon_slave_firsttransfer;
  --~read_n_to_the_ext_flash of type read to ~p1_read_n_to_the_ext_flash, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      read_n_to_the_ext_flash <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      read_n_to_the_ext_flash <= p1_read_n_to_the_ext_flash;
    end if;

  end process;

  --~p1_read_n_to_the_ext_flash assignment, which is an e_mux
  p1_read_n_to_the_ext_flash <= NOT (((((((internal_niosII_system_burst_12_downstream_granted_ext_flash_s1 AND niosII_system_burst_12_downstream_read)) OR ((internal_niosII_system_burst_13_downstream_granted_ext_flash_s1 AND niosII_system_burst_13_downstream_read)))) AND NOT tri_state_bridge_avalon_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (ext_flash_s1_wait_counter))<std_logic_vector'("00000000000000000000000000010000"))))));
  --~write_n_to_the_ext_flash of type write to ~p1_write_n_to_the_ext_flash, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      write_n_to_the_ext_flash <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      write_n_to_the_ext_flash <= p1_write_n_to_the_ext_flash;
    end if;

  end process;

  --~p1_write_n_to_the_ext_flash assignment, which is an e_mux
  p1_write_n_to_the_ext_flash <= NOT (((((((((internal_niosII_system_burst_12_downstream_granted_ext_flash_s1 AND niosII_system_burst_12_downstream_write)) OR ((internal_niosII_system_burst_13_downstream_granted_ext_flash_s1 AND niosII_system_burst_13_downstream_write)))) AND NOT tri_state_bridge_avalon_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (ext_flash_s1_wait_counter))>=std_logic_vector'("00000000000000000000000000000100"))))) AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (ext_flash_s1_wait_counter))<std_logic_vector'("00000000000000000000000000010100"))))) AND ext_flash_s1_pretend_byte_enable));
  --address_to_the_ext_flash of type address to p1_address_to_the_ext_flash, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      address_to_the_ext_flash <= std_logic_vector'("0000000000000000000000");
    elsif clk'event and clk = '1' then
      address_to_the_ext_flash <= p1_address_to_the_ext_flash;
    end if;

  end process;

  --p1_address_to_the_ext_flash mux, which is an e_mux
  p1_address_to_the_ext_flash <= A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_12_downstream_granted_ext_flash_s1)) = '1'), niosII_system_burst_12_downstream_address_to_slave, niosII_system_burst_13_downstream_address_to_slave);
  --d1_tri_state_bridge_avalon_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_tri_state_bridge_avalon_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_tri_state_bridge_avalon_slave_end_xfer <= tri_state_bridge_avalon_slave_end_xfer;
    end if;

  end process;

  --ext_flash_s1_waits_for_read in a cycle, which is an e_mux
  ext_flash_s1_waits_for_read <= ext_flash_s1_in_a_read_cycle AND wait_for_ext_flash_s1_counter;
  --ext_flash_s1_in_a_read_cycle assignment, which is an e_assign
  ext_flash_s1_in_a_read_cycle <= ((internal_niosII_system_burst_12_downstream_granted_ext_flash_s1 AND niosII_system_burst_12_downstream_read)) OR ((internal_niosII_system_burst_13_downstream_granted_ext_flash_s1 AND niosII_system_burst_13_downstream_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= ext_flash_s1_in_a_read_cycle;
  --ext_flash_s1_waits_for_write in a cycle, which is an e_mux
  ext_flash_s1_waits_for_write <= ext_flash_s1_in_a_write_cycle AND wait_for_ext_flash_s1_counter;
  --ext_flash_s1_in_a_write_cycle assignment, which is an e_assign
  ext_flash_s1_in_a_write_cycle <= ((internal_niosII_system_burst_12_downstream_granted_ext_flash_s1 AND niosII_system_burst_12_downstream_write)) OR ((internal_niosII_system_burst_13_downstream_granted_ext_flash_s1 AND niosII_system_burst_13_downstream_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= ext_flash_s1_in_a_write_cycle;
  internal_ext_flash_s1_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("000000000000000000000000000") & (ext_flash_s1_wait_counter)) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_flash_s1_wait_counter <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      ext_flash_s1_wait_counter <= ext_flash_s1_counter_load_value;
    end if;

  end process;

  ext_flash_s1_counter_load_value <= A_EXT (A_WE_StdLogicVector((std_logic'(((ext_flash_s1_in_a_read_cycle AND tri_state_bridge_avalon_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000010010"), A_WE_StdLogicVector((std_logic'(((ext_flash_s1_in_a_write_cycle AND tri_state_bridge_avalon_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000010110"), A_WE_StdLogicVector((std_logic'((NOT internal_ext_flash_s1_wait_counter_eq_0)) = '1'), ((std_logic_vector'("0000000000000000000000000000") & (ext_flash_s1_wait_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000")))), 5);
  wait_for_ext_flash_s1_counter <= tri_state_bridge_avalon_slave_begins_xfer OR NOT internal_ext_flash_s1_wait_counter_eq_0;
  --ext_flash_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  ext_flash_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_12_downstream_granted_ext_flash_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_12_downstream_byteenable))), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_13_downstream_granted_ext_flash_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_13_downstream_byteenable))), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))));
  --vhdl renameroo for output signals
  ext_flash_s1_wait_counter_eq_0 <= internal_ext_flash_s1_wait_counter_eq_0;
  --vhdl renameroo for output signals
  niosII_system_burst_12_downstream_granted_ext_flash_s1 <= internal_niosII_system_burst_12_downstream_granted_ext_flash_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 <= internal_niosII_system_burst_12_downstream_qualified_request_ext_flash_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_12_downstream_requests_ext_flash_s1 <= internal_niosII_system_burst_12_downstream_requests_ext_flash_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_13_downstream_granted_ext_flash_s1 <= internal_niosII_system_burst_13_downstream_granted_ext_flash_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 <= internal_niosII_system_burst_13_downstream_qualified_request_ext_flash_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_13_downstream_requests_ext_flash_s1 <= internal_niosII_system_burst_13_downstream_requests_ext_flash_s1;
--synthesis translate_off
    --incoming_data_to_and_from_the_ext_flash_bit_0_is_x x check, which is an e_assign_is_x
    incoming_data_to_and_from_the_ext_flash_bit_0_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_data_to_and_from_the_ext_flash(0))), '1','0');
    --Crush incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0[0] Xs to 0, which is an e_assign
    incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0(0) <= A_WE_StdLogic((std_logic'(incoming_data_to_and_from_the_ext_flash_bit_0_is_x) = '1'), std_logic'('0'), incoming_data_to_and_from_the_ext_flash(0));
    --incoming_data_to_and_from_the_ext_flash_bit_1_is_x x check, which is an e_assign_is_x
    incoming_data_to_and_from_the_ext_flash_bit_1_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_data_to_and_from_the_ext_flash(1))), '1','0');
    --Crush incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0[1] Xs to 0, which is an e_assign
    incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0(1) <= A_WE_StdLogic((std_logic'(incoming_data_to_and_from_the_ext_flash_bit_1_is_x) = '1'), std_logic'('0'), incoming_data_to_and_from_the_ext_flash(1));
    --incoming_data_to_and_from_the_ext_flash_bit_2_is_x x check, which is an e_assign_is_x
    incoming_data_to_and_from_the_ext_flash_bit_2_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_data_to_and_from_the_ext_flash(2))), '1','0');
    --Crush incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0[2] Xs to 0, which is an e_assign
    incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0(2) <= A_WE_StdLogic((std_logic'(incoming_data_to_and_from_the_ext_flash_bit_2_is_x) = '1'), std_logic'('0'), incoming_data_to_and_from_the_ext_flash(2));
    --incoming_data_to_and_from_the_ext_flash_bit_3_is_x x check, which is an e_assign_is_x
    incoming_data_to_and_from_the_ext_flash_bit_3_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_data_to_and_from_the_ext_flash(3))), '1','0');
    --Crush incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0[3] Xs to 0, which is an e_assign
    incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0(3) <= A_WE_StdLogic((std_logic'(incoming_data_to_and_from_the_ext_flash_bit_3_is_x) = '1'), std_logic'('0'), incoming_data_to_and_from_the_ext_flash(3));
    --incoming_data_to_and_from_the_ext_flash_bit_4_is_x x check, which is an e_assign_is_x
    incoming_data_to_and_from_the_ext_flash_bit_4_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_data_to_and_from_the_ext_flash(4))), '1','0');
    --Crush incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0[4] Xs to 0, which is an e_assign
    incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0(4) <= A_WE_StdLogic((std_logic'(incoming_data_to_and_from_the_ext_flash_bit_4_is_x) = '1'), std_logic'('0'), incoming_data_to_and_from_the_ext_flash(4));
    --incoming_data_to_and_from_the_ext_flash_bit_5_is_x x check, which is an e_assign_is_x
    incoming_data_to_and_from_the_ext_flash_bit_5_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_data_to_and_from_the_ext_flash(5))), '1','0');
    --Crush incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0[5] Xs to 0, which is an e_assign
    incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0(5) <= A_WE_StdLogic((std_logic'(incoming_data_to_and_from_the_ext_flash_bit_5_is_x) = '1'), std_logic'('0'), incoming_data_to_and_from_the_ext_flash(5));
    --incoming_data_to_and_from_the_ext_flash_bit_6_is_x x check, which is an e_assign_is_x
    incoming_data_to_and_from_the_ext_flash_bit_6_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_data_to_and_from_the_ext_flash(6))), '1','0');
    --Crush incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0[6] Xs to 0, which is an e_assign
    incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0(6) <= A_WE_StdLogic((std_logic'(incoming_data_to_and_from_the_ext_flash_bit_6_is_x) = '1'), std_logic'('0'), incoming_data_to_and_from_the_ext_flash(6));
    --incoming_data_to_and_from_the_ext_flash_bit_7_is_x x check, which is an e_assign_is_x
    incoming_data_to_and_from_the_ext_flash_bit_7_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_data_to_and_from_the_ext_flash(7))), '1','0');
    --Crush incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0[7] Xs to 0, which is an e_assign
    incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0(7) <= A_WE_StdLogic((std_logic'(incoming_data_to_and_from_the_ext_flash_bit_7_is_x) = '1'), std_logic'('0'), incoming_data_to_and_from_the_ext_flash(7));
    --ext_flash/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_12/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line206 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_12_downstream_requests_ext_flash_s1 AND to_std_logic((((std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_12_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line206, now);
          write(write_line206, string'(": "));
          write(write_line206, string'("niosII_system_burst_12/downstream drove 0 on its 'arbitrationshare' port while accessing slave ext_flash/s1"));
          write(output, write_line206.all);
          deallocate (write_line206);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_12/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line207 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_12_downstream_requests_ext_flash_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_12_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line207, now);
          write(write_line207, string'(": "));
          write(write_line207, string'("niosII_system_burst_12/downstream drove 0 on its 'burstcount' port while accessing slave ext_flash/s1"));
          write(output, write_line207.all);
          deallocate (write_line207);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_13/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line208 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_13_downstream_requests_ext_flash_s1 AND to_std_logic((((std_logic_vector'("00000000000000000000000000") & (niosII_system_burst_13_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line208, now);
          write(write_line208, string'(": "));
          write(write_line208, string'("niosII_system_burst_13/downstream drove 0 on its 'arbitrationshare' port while accessing slave ext_flash/s1"));
          write(output, write_line208.all);
          deallocate (write_line208);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_13/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line209 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_13_downstream_requests_ext_flash_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_13_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line209, now);
          write(write_line209, string'(": "));
          write(write_line209, string'("niosII_system_burst_13/downstream drove 0 on its 'burstcount' port while accessing slave ext_flash/s1"));
          write(output, write_line209.all);
          deallocate (write_line209);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line210 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_12_downstream_granted_ext_flash_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_13_downstream_granted_ext_flash_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line210, now);
          write(write_line210, string'(": "));
          write(write_line210, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line210.all);
          deallocate (write_line210);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line211 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(niosII_system_burst_12_downstream_saved_grant_ext_flash_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(niosII_system_burst_13_downstream_saved_grant_ext_flash_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line211, now);
          write(write_line211, string'(": "));
          write(write_line211, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line211.all);
          deallocate (write_line211);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on
--synthesis read_comments_as_HDL on
--    
--    incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 <= incoming_data_to_and_from_the_ext_flash;
--synthesis read_comments_as_HDL off

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tri_state_bridge_bridge_arbitrator is 
end entity tri_state_bridge_bridge_arbitrator;


architecture europa of tri_state_bridge_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity tsb_avalon_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_address_to_slave : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_19_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_address_to_slave : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_20_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_system_burst_20_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_20_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_20_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_tsb_avalon_slave_end_xfer : OUT STD_LOGIC;
                 signal incoming_sram_IF_0_tsb_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_system_burst_19_downstream_granted_sram_IF_0_tsb : OUT STD_LOGIC;
                 signal niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb : OUT STD_LOGIC;
                 signal niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb : OUT STD_LOGIC;
                 signal niosII_system_burst_19_downstream_requests_sram_IF_0_tsb : OUT STD_LOGIC;
                 signal niosII_system_burst_20_downstream_granted_sram_IF_0_tsb : OUT STD_LOGIC;
                 signal niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb : OUT STD_LOGIC;
                 signal niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb : OUT STD_LOGIC;
                 signal niosII_system_burst_20_downstream_requests_sram_IF_0_tsb : OUT STD_LOGIC;
                 signal sram_IF_0_tsb_address : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal sram_IF_0_tsb_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sram_IF_0_tsb_chipselect_n : OUT STD_LOGIC;
                 signal sram_IF_0_tsb_data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sram_IF_0_tsb_outputenable_n : OUT STD_LOGIC;
                 signal sram_IF_0_tsb_write_n : OUT STD_LOGIC
              );
end entity tsb_avalon_slave_arbitrator;


architecture europa of tsb_avalon_slave_arbitrator is
                signal d1_in_a_write_cycle :  STD_LOGIC;
                signal d1_outgoing_sram_IF_0_tsb_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_tsb_avalon_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb :  STD_LOGIC;
                signal internal_niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb :  STD_LOGIC;
                signal internal_niosII_system_burst_19_downstream_requests_sram_IF_0_tsb :  STD_LOGIC;
                signal internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb :  STD_LOGIC;
                signal internal_niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb :  STD_LOGIC;
                signal internal_niosII_system_burst_20_downstream_requests_sram_IF_0_tsb :  STD_LOGIC;
                signal last_cycle_niosII_system_burst_19_downstream_granted_slave_sram_IF_0_tsb :  STD_LOGIC;
                signal last_cycle_niosII_system_burst_20_downstream_granted_slave_sram_IF_0_tsb :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register_in :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_saved_grant_sram_IF_0_tsb :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register_in :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_saved_grant_sram_IF_0_tsb :  STD_LOGIC;
                signal outgoing_sram_IF_0_tsb_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_sram_IF_0_tsb_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal p1_sram_IF_0_tsb_byteenable_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_sram_IF_0_tsb_chipselect_n :  STD_LOGIC;
                signal p1_sram_IF_0_tsb_outputenable_n :  STD_LOGIC;
                signal p1_sram_IF_0_tsb_write_n :  STD_LOGIC;
                signal sram_IF_0_tsb_in_a_read_cycle :  STD_LOGIC;
                signal sram_IF_0_tsb_in_a_write_cycle :  STD_LOGIC;
                signal sram_IF_0_tsb_waits_for_read :  STD_LOGIC;
                signal sram_IF_0_tsb_waits_for_write :  STD_LOGIC;
                signal sram_IF_0_tsb_with_write_latency :  STD_LOGIC;
                signal time_to_write :  STD_LOGIC;
                signal tsb_avalon_slave_allgrants :  STD_LOGIC;
                signal tsb_avalon_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal tsb_avalon_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal tsb_avalon_slave_any_continuerequest :  STD_LOGIC;
                signal tsb_avalon_slave_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tsb_avalon_slave_arb_counter_enable :  STD_LOGIC;
                signal tsb_avalon_slave_arb_share_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal tsb_avalon_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal tsb_avalon_slave_arb_share_set_values :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal tsb_avalon_slave_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tsb_avalon_slave_arbitration_holdoff_internal :  STD_LOGIC;
                signal tsb_avalon_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal tsb_avalon_slave_begins_xfer :  STD_LOGIC;
                signal tsb_avalon_slave_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tsb_avalon_slave_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tsb_avalon_slave_end_xfer :  STD_LOGIC;
                signal tsb_avalon_slave_firsttransfer :  STD_LOGIC;
                signal tsb_avalon_slave_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tsb_avalon_slave_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tsb_avalon_slave_non_bursting_master_requests :  STD_LOGIC;
                signal tsb_avalon_slave_read_pending :  STD_LOGIC;
                signal tsb_avalon_slave_reg_firsttransfer :  STD_LOGIC;
                signal tsb_avalon_slave_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tsb_avalon_slave_slavearbiterlockenable :  STD_LOGIC;
                signal tsb_avalon_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal tsb_avalon_slave_unreg_firsttransfer :  STD_LOGIC;
                signal tsb_avalon_slave_write_pending :  STD_LOGIC;
                signal wait_for_sram_IF_0_tsb_counter :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of d1_in_a_write_cycle : signal is "FAST_OUTPUT_ENABLE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of d1_outgoing_sram_IF_0_tsb_data : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of incoming_sram_IF_0_tsb_data : signal is "FAST_INPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of sram_IF_0_tsb_address : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of sram_IF_0_tsb_byteenable_n : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of sram_IF_0_tsb_chipselect_n : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of sram_IF_0_tsb_outputenable_n : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of sram_IF_0_tsb_write_n : signal is "FAST_OUTPUT_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT tsb_avalon_slave_end_xfer;
    end if;

  end process;

  tsb_avalon_slave_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb OR internal_niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb));
  internal_niosII_system_burst_19_downstream_requests_sram_IF_0_tsb <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_19_downstream_read OR niosII_system_burst_19_downstream_write)))))));
  --~sram_IF_0_tsb_chipselect_n of type chipselect to ~p1_sram_IF_0_tsb_chipselect_n, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sram_IF_0_tsb_chipselect_n <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      sram_IF_0_tsb_chipselect_n <= p1_sram_IF_0_tsb_chipselect_n;
    end if;

  end process;

  tsb_avalon_slave_write_pending <= std_logic'('0');
  --tsb/avalon_slave read pending calc, which is an e_assign
  tsb_avalon_slave_read_pending <= std_logic'('0');
  --tsb_avalon_slave_arb_share_counter set values, which is an e_mux
  tsb_avalon_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_19_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_20_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_19_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_20_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001"))))), 5);
  --tsb_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  tsb_avalon_slave_non_bursting_master_requests <= std_logic'('0');
  --tsb_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  tsb_avalon_slave_any_bursting_master_saved_grant <= ((niosII_system_burst_19_downstream_saved_grant_sram_IF_0_tsb OR niosII_system_burst_20_downstream_saved_grant_sram_IF_0_tsb) OR niosII_system_burst_19_downstream_saved_grant_sram_IF_0_tsb) OR niosII_system_burst_20_downstream_saved_grant_sram_IF_0_tsb;
  --tsb_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  tsb_avalon_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(tsb_avalon_slave_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (tsb_avalon_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(tsb_avalon_slave_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (tsb_avalon_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 5);
  --tsb_avalon_slave_allgrants all slave grants, which is an e_mux
  tsb_avalon_slave_allgrants <= (((or_reduce(tsb_avalon_slave_grant_vector)) OR (or_reduce(tsb_avalon_slave_grant_vector))) OR (or_reduce(tsb_avalon_slave_grant_vector))) OR (or_reduce(tsb_avalon_slave_grant_vector));
  --tsb_avalon_slave_end_xfer assignment, which is an e_assign
  tsb_avalon_slave_end_xfer <= NOT ((sram_IF_0_tsb_waits_for_read OR sram_IF_0_tsb_waits_for_write));
  --end_xfer_arb_share_counter_term_tsb_avalon_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_tsb_avalon_slave <= tsb_avalon_slave_end_xfer AND (((NOT tsb_avalon_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --tsb_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  tsb_avalon_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_tsb_avalon_slave AND tsb_avalon_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_tsb_avalon_slave AND NOT tsb_avalon_slave_non_bursting_master_requests));
  --tsb_avalon_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tsb_avalon_slave_arb_share_counter <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(tsb_avalon_slave_arb_counter_enable) = '1' then 
        tsb_avalon_slave_arb_share_counter <= tsb_avalon_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --tsb_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tsb_avalon_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(tsb_avalon_slave_master_qreq_vector) AND end_xfer_arb_share_counter_term_tsb_avalon_slave)) OR ((end_xfer_arb_share_counter_term_tsb_avalon_slave AND NOT tsb_avalon_slave_non_bursting_master_requests)))) = '1' then 
        tsb_avalon_slave_slavearbiterlockenable <= or_reduce(tsb_avalon_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_19/downstream tsb/avalon_slave arbiterlock, which is an e_assign
  niosII_system_burst_19_downstream_arbiterlock <= tsb_avalon_slave_slavearbiterlockenable AND niosII_system_burst_19_downstream_continuerequest;
  --tsb_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  tsb_avalon_slave_slavearbiterlockenable2 <= or_reduce(tsb_avalon_slave_arb_share_counter_next_value);
  --niosII_system_burst_19/downstream tsb/avalon_slave arbiterlock2, which is an e_assign
  niosII_system_burst_19_downstream_arbiterlock2 <= tsb_avalon_slave_slavearbiterlockenable2 AND niosII_system_burst_19_downstream_continuerequest;
  --niosII_system_burst_20/downstream tsb/avalon_slave arbiterlock, which is an e_assign
  niosII_system_burst_20_downstream_arbiterlock <= tsb_avalon_slave_slavearbiterlockenable AND niosII_system_burst_20_downstream_continuerequest;
  --niosII_system_burst_20/downstream tsb/avalon_slave arbiterlock2, which is an e_assign
  niosII_system_burst_20_downstream_arbiterlock2 <= tsb_avalon_slave_slavearbiterlockenable2 AND niosII_system_burst_20_downstream_continuerequest;
  --niosII_system_burst_20/downstream granted sram_IF_0/tsb last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_niosII_system_burst_20_downstream_granted_slave_sram_IF_0_tsb <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_niosII_system_burst_20_downstream_granted_slave_sram_IF_0_tsb <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(niosII_system_burst_20_downstream_saved_grant_sram_IF_0_tsb) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tsb_avalon_slave_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_20_downstream_granted_slave_sram_IF_0_tsb))))));
    end if;

  end process;

  --niosII_system_burst_20_downstream_continuerequest continued request, which is an e_mux
  niosII_system_burst_20_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_20_downstream_granted_slave_sram_IF_0_tsb))) AND std_logic_vector'("00000000000000000000000000000001")));
  --tsb_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  tsb_avalon_slave_any_continuerequest <= niosII_system_burst_20_downstream_continuerequest OR niosII_system_burst_19_downstream_continuerequest;
  internal_niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb <= internal_niosII_system_burst_19_downstream_requests_sram_IF_0_tsb AND NOT (((((niosII_system_burst_19_downstream_read AND ((tsb_avalon_slave_write_pending OR (tsb_avalon_slave_read_pending))))) OR (((tsb_avalon_slave_read_pending) AND niosII_system_burst_19_downstream_write))) OR niosII_system_burst_20_downstream_arbiterlock));
  --niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register_in mux for readlatency shift register, which is an e_mux
  niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register_in <= (internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb AND niosII_system_burst_19_downstream_read) AND NOT sram_IF_0_tsb_waits_for_read;
  --shift register p1 niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register <= A_EXT ((niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register & A_ToStdLogicVector(niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register_in)), 2);
  --niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register <= p1_niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register;
    end if;

  end process;

  --local readdatavalid niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb, which is an e_mux
  niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb <= niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb_shift_register(1);
  --sram_IF_0_tsb_data register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      incoming_sram_IF_0_tsb_data <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      incoming_sram_IF_0_tsb_data <= sram_IF_0_tsb_data;
    end if;

  end process;

  --sram_IF_0_tsb_with_write_latency assignment, which is an e_assign
  sram_IF_0_tsb_with_write_latency <= in_a_write_cycle AND ((internal_niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb OR internal_niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb));
  --time to write the data, which is an e_mux
  time_to_write <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((sram_IF_0_tsb_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((sram_IF_0_tsb_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), std_logic_vector'("00000000000000000000000000000000"))));
  --d1_outgoing_sram_IF_0_tsb_data register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_outgoing_sram_IF_0_tsb_data <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      d1_outgoing_sram_IF_0_tsb_data <= outgoing_sram_IF_0_tsb_data;
    end if;

  end process;

  --write cycle delayed by 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_in_a_write_cycle <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_in_a_write_cycle <= time_to_write;
    end if;

  end process;

  --d1_outgoing_sram_IF_0_tsb_data tristate driver, which is an e_assign
  sram_IF_0_tsb_data <= A_WE_StdLogicVector((std_logic'((d1_in_a_write_cycle)) = '1'), d1_outgoing_sram_IF_0_tsb_data, A_REP(std_logic'('Z'), 16));
  --outgoing_sram_IF_0_tsb_data mux, which is an e_mux
  outgoing_sram_IF_0_tsb_data <= A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb)) = '1'), niosII_system_burst_19_downstream_writedata, niosII_system_burst_20_downstream_writedata);
  internal_niosII_system_burst_20_downstream_requests_sram_IF_0_tsb <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_20_downstream_read OR niosII_system_burst_20_downstream_write)))))));
  --niosII_system_burst_19/downstream granted sram_IF_0/tsb last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_niosII_system_burst_19_downstream_granted_slave_sram_IF_0_tsb <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_niosII_system_burst_19_downstream_granted_slave_sram_IF_0_tsb <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(niosII_system_burst_19_downstream_saved_grant_sram_IF_0_tsb) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tsb_avalon_slave_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_19_downstream_granted_slave_sram_IF_0_tsb))))));
    end if;

  end process;

  --niosII_system_burst_19_downstream_continuerequest continued request, which is an e_mux
  niosII_system_burst_19_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_niosII_system_burst_19_downstream_granted_slave_sram_IF_0_tsb))) AND std_logic_vector'("00000000000000000000000000000001")));
  internal_niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb <= internal_niosII_system_burst_20_downstream_requests_sram_IF_0_tsb AND NOT (((((niosII_system_burst_20_downstream_read AND ((tsb_avalon_slave_write_pending OR (tsb_avalon_slave_read_pending))))) OR (((tsb_avalon_slave_read_pending) AND niosII_system_burst_20_downstream_write))) OR niosII_system_burst_19_downstream_arbiterlock));
  --niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register_in mux for readlatency shift register, which is an e_mux
  niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register_in <= (internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb AND niosII_system_burst_20_downstream_read) AND NOT sram_IF_0_tsb_waits_for_read;
  --shift register p1 niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register <= A_EXT ((niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register & A_ToStdLogicVector(niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register_in)), 2);
  --niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register <= p1_niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register;
    end if;

  end process;

  --local readdatavalid niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb, which is an e_mux
  niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb <= niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb_shift_register(1);
  --allow new arb cycle for tsb/avalon_slave, which is an e_assign
  tsb_avalon_slave_allow_new_arb_cycle <= NOT niosII_system_burst_19_downstream_arbiterlock AND NOT niosII_system_burst_20_downstream_arbiterlock;
  --niosII_system_burst_20/downstream assignment into master qualified-requests vector for sram_IF_0/tsb, which is an e_assign
  tsb_avalon_slave_master_qreq_vector(0) <= internal_niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb;
  --niosII_system_burst_20/downstream grant sram_IF_0/tsb, which is an e_assign
  internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb <= tsb_avalon_slave_grant_vector(0);
  --niosII_system_burst_20/downstream saved-grant sram_IF_0/tsb, which is an e_assign
  niosII_system_burst_20_downstream_saved_grant_sram_IF_0_tsb <= tsb_avalon_slave_arb_winner(0);
  --niosII_system_burst_19/downstream assignment into master qualified-requests vector for sram_IF_0/tsb, which is an e_assign
  tsb_avalon_slave_master_qreq_vector(1) <= internal_niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb;
  --niosII_system_burst_19/downstream grant sram_IF_0/tsb, which is an e_assign
  internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb <= tsb_avalon_slave_grant_vector(1);
  --niosII_system_burst_19/downstream saved-grant sram_IF_0/tsb, which is an e_assign
  niosII_system_burst_19_downstream_saved_grant_sram_IF_0_tsb <= tsb_avalon_slave_arb_winner(1);
  --tsb/avalon_slave chosen-master double-vector, which is an e_assign
  tsb_avalon_slave_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((tsb_avalon_slave_master_qreq_vector & tsb_avalon_slave_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT tsb_avalon_slave_master_qreq_vector & NOT tsb_avalon_slave_master_qreq_vector))) + (std_logic_vector'("000") & (tsb_avalon_slave_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  tsb_avalon_slave_arb_winner <= A_WE_StdLogicVector((std_logic'(((tsb_avalon_slave_allow_new_arb_cycle AND or_reduce(tsb_avalon_slave_grant_vector)))) = '1'), tsb_avalon_slave_grant_vector, tsb_avalon_slave_saved_chosen_master_vector);
  --saved tsb_avalon_slave_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tsb_avalon_slave_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(tsb_avalon_slave_allow_new_arb_cycle) = '1' then 
        tsb_avalon_slave_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(tsb_avalon_slave_grant_vector)) = '1'), tsb_avalon_slave_grant_vector, tsb_avalon_slave_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  tsb_avalon_slave_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((tsb_avalon_slave_chosen_master_double_vector(1) OR tsb_avalon_slave_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((tsb_avalon_slave_chosen_master_double_vector(0) OR tsb_avalon_slave_chosen_master_double_vector(2)))));
  --tsb/avalon_slave chosen master rotated left, which is an e_assign
  tsb_avalon_slave_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(tsb_avalon_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(tsb_avalon_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --tsb/avalon_slave's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tsb_avalon_slave_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(tsb_avalon_slave_grant_vector)) = '1' then 
        tsb_avalon_slave_arb_addend <= A_WE_StdLogicVector((std_logic'(tsb_avalon_slave_end_xfer) = '1'), tsb_avalon_slave_chosen_master_rot_left, tsb_avalon_slave_grant_vector);
      end if;
    end if;

  end process;

  --~sram_IF_0_tsb_outputenable_n of type outputenable to ~p1_sram_IF_0_tsb_outputenable_n, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sram_IF_0_tsb_outputenable_n <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      sram_IF_0_tsb_outputenable_n <= p1_sram_IF_0_tsb_outputenable_n;
    end if;

  end process;

  --~p1_sram_IF_0_tsb_outputenable_n assignment, which is an e_mux
  p1_sram_IF_0_tsb_outputenable_n <= NOT sram_IF_0_tsb_in_a_read_cycle;
  p1_sram_IF_0_tsb_chipselect_n <= NOT ((internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb OR internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb));
  --tsb_avalon_slave_firsttransfer first transaction, which is an e_assign
  tsb_avalon_slave_firsttransfer <= A_WE_StdLogic((std_logic'(tsb_avalon_slave_begins_xfer) = '1'), tsb_avalon_slave_unreg_firsttransfer, tsb_avalon_slave_reg_firsttransfer);
  --tsb_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  tsb_avalon_slave_unreg_firsttransfer <= NOT ((tsb_avalon_slave_slavearbiterlockenable AND tsb_avalon_slave_any_continuerequest));
  --tsb_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tsb_avalon_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(tsb_avalon_slave_begins_xfer) = '1' then 
        tsb_avalon_slave_reg_firsttransfer <= tsb_avalon_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --tsb_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  tsb_avalon_slave_beginbursttransfer_internal <= tsb_avalon_slave_begins_xfer;
  --tsb_avalon_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  tsb_avalon_slave_arbitration_holdoff_internal <= tsb_avalon_slave_begins_xfer AND tsb_avalon_slave_firsttransfer;
  --~sram_IF_0_tsb_write_n of type write to ~p1_sram_IF_0_tsb_write_n, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sram_IF_0_tsb_write_n <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      sram_IF_0_tsb_write_n <= p1_sram_IF_0_tsb_write_n;
    end if;

  end process;

  --~sram_IF_0_tsb_byteenable_n of type byteenable to ~p1_sram_IF_0_tsb_byteenable_n, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sram_IF_0_tsb_byteenable_n <= A_EXT (NOT std_logic_vector'("00000000000000000000000000000000"), 2);
    elsif clk'event and clk = '1' then
      sram_IF_0_tsb_byteenable_n <= p1_sram_IF_0_tsb_byteenable_n;
    end if;

  end process;

  --~p1_sram_IF_0_tsb_write_n assignment, which is an e_mux
  p1_sram_IF_0_tsb_write_n <= NOT ((((internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb AND niosII_system_burst_19_downstream_write)) OR ((internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb AND niosII_system_burst_20_downstream_write))));
  --sram_IF_0_tsb_address of type address to p1_sram_IF_0_tsb_address, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sram_IF_0_tsb_address <= std_logic_vector'("0000000000000000000");
    elsif clk'event and clk = '1' then
      sram_IF_0_tsb_address <= p1_sram_IF_0_tsb_address;
    end if;

  end process;

  --p1_sram_IF_0_tsb_address mux, which is an e_mux
  p1_sram_IF_0_tsb_address <= A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb)) = '1'), niosII_system_burst_19_downstream_address_to_slave, niosII_system_burst_20_downstream_address_to_slave);
  --d1_tsb_avalon_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_tsb_avalon_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_tsb_avalon_slave_end_xfer <= tsb_avalon_slave_end_xfer;
    end if;

  end process;

  --sram_IF_0_tsb_waits_for_read in a cycle, which is an e_mux
  sram_IF_0_tsb_waits_for_read <= sram_IF_0_tsb_in_a_read_cycle AND tsb_avalon_slave_begins_xfer;
  --sram_IF_0_tsb_in_a_read_cycle assignment, which is an e_assign
  sram_IF_0_tsb_in_a_read_cycle <= ((internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb AND niosII_system_burst_19_downstream_read)) OR ((internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb AND niosII_system_burst_20_downstream_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sram_IF_0_tsb_in_a_read_cycle;
  --sram_IF_0_tsb_waits_for_write in a cycle, which is an e_mux
  sram_IF_0_tsb_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sram_IF_0_tsb_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sram_IF_0_tsb_in_a_write_cycle assignment, which is an e_assign
  sram_IF_0_tsb_in_a_write_cycle <= ((internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb AND niosII_system_burst_19_downstream_write)) OR ((internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb AND niosII_system_burst_20_downstream_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sram_IF_0_tsb_in_a_write_cycle;
  wait_for_sram_IF_0_tsb_counter <= std_logic'('0');
  --~p1_sram_IF_0_tsb_byteenable_n byte enable port mux, which is an e_mux
  p1_sram_IF_0_tsb_byteenable_n <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_19_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (niosII_system_burst_20_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))))), 2);
  --vhdl renameroo for output signals
  niosII_system_burst_19_downstream_granted_sram_IF_0_tsb <= internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb;
  --vhdl renameroo for output signals
  niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb <= internal_niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb;
  --vhdl renameroo for output signals
  niosII_system_burst_19_downstream_requests_sram_IF_0_tsb <= internal_niosII_system_burst_19_downstream_requests_sram_IF_0_tsb;
  --vhdl renameroo for output signals
  niosII_system_burst_20_downstream_granted_sram_IF_0_tsb <= internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb;
  --vhdl renameroo for output signals
  niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb <= internal_niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb;
  --vhdl renameroo for output signals
  niosII_system_burst_20_downstream_requests_sram_IF_0_tsb <= internal_niosII_system_burst_20_downstream_requests_sram_IF_0_tsb;
--synthesis translate_off
    --sram_IF_0/tsb enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_19/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line212 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_19_downstream_requests_sram_IF_0_tsb AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_19_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line212, now);
          write(write_line212, string'(": "));
          write(write_line212, string'("niosII_system_burst_19/downstream drove 0 on its 'arbitrationshare' port while accessing slave sram_IF_0/tsb"));
          write(output, write_line212.all);
          deallocate (write_line212);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_19/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line213 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_19_downstream_requests_sram_IF_0_tsb AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_19_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line213, now);
          write(write_line213, string'(": "));
          write(write_line213, string'("niosII_system_burst_19/downstream drove 0 on its 'burstcount' port while accessing slave sram_IF_0/tsb"));
          write(output, write_line213.all);
          deallocate (write_line213);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_20/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line214 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_20_downstream_requests_sram_IF_0_tsb AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_20_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line214, now);
          write(write_line214, string'(": "));
          write(write_line214, string'("niosII_system_burst_20/downstream drove 0 on its 'arbitrationshare' port while accessing slave sram_IF_0/tsb"));
          write(output, write_line214.all);
          deallocate (write_line214);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_20/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line215 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_20_downstream_requests_sram_IF_0_tsb AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_20_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line215, now);
          write(write_line215, string'(": "));
          write(write_line215, string'("niosII_system_burst_20/downstream drove 0 on its 'burstcount' port while accessing slave sram_IF_0/tsb"));
          write(output, write_line215.all);
          deallocate (write_line215);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line216 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_19_downstream_granted_sram_IF_0_tsb))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_niosII_system_burst_20_downstream_granted_sram_IF_0_tsb))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line216, now);
          write(write_line216, string'(": "));
          write(write_line216, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line216.all);
          deallocate (write_line216);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line217 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(niosII_system_burst_19_downstream_saved_grant_sram_IF_0_tsb))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(niosII_system_burst_20_downstream_saved_grant_sram_IF_0_tsb))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line217, now);
          write(write_line217, string'(": "));
          write(write_line217, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line217.all);
          deallocate (write_line217);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tsb_bridge_arbitrator is 
end entity tsb_bridge_arbitrator;


architecture europa of tsb_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity uart_0_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_17_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_17_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_17_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_17_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal uart_0_s1_dataavailable : IN STD_LOGIC;
                 signal uart_0_s1_irq : IN STD_LOGIC;
                 signal uart_0_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal uart_0_s1_readyfordata : IN STD_LOGIC;

              -- outputs:
                 signal d1_uart_0_s1_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_17_downstream_granted_uart_0_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_17_downstream_qualified_request_uart_0_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_17_downstream_read_data_valid_uart_0_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_17_downstream_requests_uart_0_s1 : OUT STD_LOGIC;
                 signal uart_0_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal uart_0_s1_begintransfer : OUT STD_LOGIC;
                 signal uart_0_s1_chipselect : OUT STD_LOGIC;
                 signal uart_0_s1_dataavailable_from_sa : OUT STD_LOGIC;
                 signal uart_0_s1_irq_from_sa : OUT STD_LOGIC;
                 signal uart_0_s1_read_n : OUT STD_LOGIC;
                 signal uart_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal uart_0_s1_readyfordata_from_sa : OUT STD_LOGIC;
                 signal uart_0_s1_reset_n : OUT STD_LOGIC;
                 signal uart_0_s1_write_n : OUT STD_LOGIC;
                 signal uart_0_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity uart_0_s1_arbitrator;


architecture europa of uart_0_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_uart_0_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_17_downstream_granted_uart_0_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_17_downstream_qualified_request_uart_0_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_17_downstream_requests_uart_0_s1 :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_saved_grant_uart_0_s1 :  STD_LOGIC;
                signal uart_0_s1_allgrants :  STD_LOGIC;
                signal uart_0_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal uart_0_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal uart_0_s1_any_continuerequest :  STD_LOGIC;
                signal uart_0_s1_arb_counter_enable :  STD_LOGIC;
                signal uart_0_s1_arb_share_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal uart_0_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal uart_0_s1_arb_share_set_values :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal uart_0_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal uart_0_s1_begins_xfer :  STD_LOGIC;
                signal uart_0_s1_end_xfer :  STD_LOGIC;
                signal uart_0_s1_firsttransfer :  STD_LOGIC;
                signal uart_0_s1_grant_vector :  STD_LOGIC;
                signal uart_0_s1_in_a_read_cycle :  STD_LOGIC;
                signal uart_0_s1_in_a_write_cycle :  STD_LOGIC;
                signal uart_0_s1_master_qreq_vector :  STD_LOGIC;
                signal uart_0_s1_non_bursting_master_requests :  STD_LOGIC;
                signal uart_0_s1_reg_firsttransfer :  STD_LOGIC;
                signal uart_0_s1_slavearbiterlockenable :  STD_LOGIC;
                signal uart_0_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal uart_0_s1_unreg_firsttransfer :  STD_LOGIC;
                signal uart_0_s1_waits_for_read :  STD_LOGIC;
                signal uart_0_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_uart_0_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT uart_0_s1_end_xfer;
    end if;

  end process;

  uart_0_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_17_downstream_qualified_request_uart_0_s1);
  --assign uart_0_s1_readdata_from_sa = uart_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart_0_s1_readdata_from_sa <= uart_0_s1_readdata;
  internal_niosII_system_burst_17_downstream_requests_uart_0_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_17_downstream_read OR niosII_system_burst_17_downstream_write)))))));
  --assign uart_0_s1_dataavailable_from_sa = uart_0_s1_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart_0_s1_dataavailable_from_sa <= uart_0_s1_dataavailable;
  --assign uart_0_s1_readyfordata_from_sa = uart_0_s1_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart_0_s1_readyfordata_from_sa <= uart_0_s1_readyfordata;
  --uart_0_s1_arb_share_counter set values, which is an e_mux
  uart_0_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_17_downstream_granted_uart_0_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_17_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --uart_0_s1_non_bursting_master_requests mux, which is an e_mux
  uart_0_s1_non_bursting_master_requests <= std_logic'('0');
  --uart_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  uart_0_s1_any_bursting_master_saved_grant <= niosII_system_burst_17_downstream_saved_grant_uart_0_s1;
  --uart_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  uart_0_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(uart_0_s1_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (uart_0_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(uart_0_s1_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (uart_0_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 5);
  --uart_0_s1_allgrants all slave grants, which is an e_mux
  uart_0_s1_allgrants <= uart_0_s1_grant_vector;
  --uart_0_s1_end_xfer assignment, which is an e_assign
  uart_0_s1_end_xfer <= NOT ((uart_0_s1_waits_for_read OR uart_0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_uart_0_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_uart_0_s1 <= uart_0_s1_end_xfer AND (((NOT uart_0_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --uart_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  uart_0_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_uart_0_s1 AND uart_0_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_uart_0_s1 AND NOT uart_0_s1_non_bursting_master_requests));
  --uart_0_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      uart_0_s1_arb_share_counter <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(uart_0_s1_arb_counter_enable) = '1' then 
        uart_0_s1_arb_share_counter <= uart_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --uart_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      uart_0_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((uart_0_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_uart_0_s1)) OR ((end_xfer_arb_share_counter_term_uart_0_s1 AND NOT uart_0_s1_non_bursting_master_requests)))) = '1' then 
        uart_0_s1_slavearbiterlockenable <= or_reduce(uart_0_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_17/downstream uart_0/s1 arbiterlock, which is an e_assign
  niosII_system_burst_17_downstream_arbiterlock <= uart_0_s1_slavearbiterlockenable AND niosII_system_burst_17_downstream_continuerequest;
  --uart_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  uart_0_s1_slavearbiterlockenable2 <= or_reduce(uart_0_s1_arb_share_counter_next_value);
  --niosII_system_burst_17/downstream uart_0/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_17_downstream_arbiterlock2 <= uart_0_s1_slavearbiterlockenable2 AND niosII_system_burst_17_downstream_continuerequest;
  --uart_0_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  uart_0_s1_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_17_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_17_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_17_downstream_qualified_request_uart_0_s1 <= internal_niosII_system_burst_17_downstream_requests_uart_0_s1 AND NOT ((niosII_system_burst_17_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_17_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_17_downstream_read_data_valid_uart_0_s1, which is an e_mux
  niosII_system_burst_17_downstream_read_data_valid_uart_0_s1 <= (internal_niosII_system_burst_17_downstream_granted_uart_0_s1 AND niosII_system_burst_17_downstream_read) AND NOT uart_0_s1_waits_for_read;
  --uart_0_s1_writedata mux, which is an e_mux
  uart_0_s1_writedata <= niosII_system_burst_17_downstream_writedata;
  --master is always granted when requested
  internal_niosII_system_burst_17_downstream_granted_uart_0_s1 <= internal_niosII_system_burst_17_downstream_qualified_request_uart_0_s1;
  --niosII_system_burst_17/downstream saved-grant uart_0/s1, which is an e_assign
  niosII_system_burst_17_downstream_saved_grant_uart_0_s1 <= internal_niosII_system_burst_17_downstream_requests_uart_0_s1;
  --allow new arb cycle for uart_0/s1, which is an e_assign
  uart_0_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  uart_0_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  uart_0_s1_master_qreq_vector <= std_logic'('1');
  uart_0_s1_begintransfer <= uart_0_s1_begins_xfer;
  --uart_0_s1_reset_n assignment, which is an e_assign
  uart_0_s1_reset_n <= reset_n;
  uart_0_s1_chipselect <= internal_niosII_system_burst_17_downstream_granted_uart_0_s1;
  --uart_0_s1_firsttransfer first transaction, which is an e_assign
  uart_0_s1_firsttransfer <= A_WE_StdLogic((std_logic'(uart_0_s1_begins_xfer) = '1'), uart_0_s1_unreg_firsttransfer, uart_0_s1_reg_firsttransfer);
  --uart_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  uart_0_s1_unreg_firsttransfer <= NOT ((uart_0_s1_slavearbiterlockenable AND uart_0_s1_any_continuerequest));
  --uart_0_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      uart_0_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(uart_0_s1_begins_xfer) = '1' then 
        uart_0_s1_reg_firsttransfer <= uart_0_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --uart_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  uart_0_s1_beginbursttransfer_internal <= uart_0_s1_begins_xfer;
  --~uart_0_s1_read_n assignment, which is an e_mux
  uart_0_s1_read_n <= NOT ((internal_niosII_system_burst_17_downstream_granted_uart_0_s1 AND niosII_system_burst_17_downstream_read));
  --~uart_0_s1_write_n assignment, which is an e_mux
  uart_0_s1_write_n <= NOT ((internal_niosII_system_burst_17_downstream_granted_uart_0_s1 AND niosII_system_burst_17_downstream_write));
  --uart_0_s1_address mux, which is an e_mux
  uart_0_s1_address <= niosII_system_burst_17_downstream_nativeaddress (2 DOWNTO 0);
  --d1_uart_0_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_uart_0_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_uart_0_s1_end_xfer <= uart_0_s1_end_xfer;
    end if;

  end process;

  --uart_0_s1_waits_for_read in a cycle, which is an e_mux
  uart_0_s1_waits_for_read <= uart_0_s1_in_a_read_cycle AND uart_0_s1_begins_xfer;
  --uart_0_s1_in_a_read_cycle assignment, which is an e_assign
  uart_0_s1_in_a_read_cycle <= internal_niosII_system_burst_17_downstream_granted_uart_0_s1 AND niosII_system_burst_17_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= uart_0_s1_in_a_read_cycle;
  --uart_0_s1_waits_for_write in a cycle, which is an e_mux
  uart_0_s1_waits_for_write <= uart_0_s1_in_a_write_cycle AND uart_0_s1_begins_xfer;
  --uart_0_s1_in_a_write_cycle assignment, which is an e_assign
  uart_0_s1_in_a_write_cycle <= internal_niosII_system_burst_17_downstream_granted_uart_0_s1 AND niosII_system_burst_17_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= uart_0_s1_in_a_write_cycle;
  wait_for_uart_0_s1_counter <= std_logic'('0');
  --assign uart_0_s1_irq_from_sa = uart_0_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart_0_s1_irq_from_sa <= uart_0_s1_irq;
  --vhdl renameroo for output signals
  niosII_system_burst_17_downstream_granted_uart_0_s1 <= internal_niosII_system_burst_17_downstream_granted_uart_0_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_17_downstream_qualified_request_uart_0_s1 <= internal_niosII_system_burst_17_downstream_qualified_request_uart_0_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_17_downstream_requests_uart_0_s1 <= internal_niosII_system_burst_17_downstream_requests_uart_0_s1;
--synthesis translate_off
    --uart_0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_17/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line218 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_17_downstream_requests_uart_0_s1 AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_17_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line218, now);
          write(write_line218, string'(": "));
          write(write_line218, string'("niosII_system_burst_17/downstream drove 0 on its 'arbitrationshare' port while accessing slave uart_0/s1"));
          write(output, write_line218.all);
          deallocate (write_line218);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_17/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line219 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_17_downstream_requests_uart_0_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_17_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line219, now);
          write(write_line219, string'(": "));
          write(write_line219, string'("niosII_system_burst_17/downstream drove 0 on its 'burstcount' port while accessing slave uart_0/s1"));
          write(output, write_line219.all);
          deallocate (write_line219);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity uart_1_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_18_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal niosII_system_burst_18_downstream_burstcount : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_latency_counter : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_system_burst_18_downstream_read : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_write : IN STD_LOGIC;
                 signal niosII_system_burst_18_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal uart_1_s1_dataavailable : IN STD_LOGIC;
                 signal uart_1_s1_irq : IN STD_LOGIC;
                 signal uart_1_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal uart_1_s1_readyfordata : IN STD_LOGIC;

              -- outputs:
                 signal d1_uart_1_s1_end_xfer : OUT STD_LOGIC;
                 signal niosII_system_burst_18_downstream_granted_uart_1_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_18_downstream_qualified_request_uart_1_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_18_downstream_read_data_valid_uart_1_s1 : OUT STD_LOGIC;
                 signal niosII_system_burst_18_downstream_requests_uart_1_s1 : OUT STD_LOGIC;
                 signal uart_1_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal uart_1_s1_begintransfer : OUT STD_LOGIC;
                 signal uart_1_s1_chipselect : OUT STD_LOGIC;
                 signal uart_1_s1_dataavailable_from_sa : OUT STD_LOGIC;
                 signal uart_1_s1_irq_from_sa : OUT STD_LOGIC;
                 signal uart_1_s1_read_n : OUT STD_LOGIC;
                 signal uart_1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal uart_1_s1_readyfordata_from_sa : OUT STD_LOGIC;
                 signal uart_1_s1_reset_n : OUT STD_LOGIC;
                 signal uart_1_s1_write_n : OUT STD_LOGIC;
                 signal uart_1_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity uart_1_s1_arbitrator;


architecture europa of uart_1_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_uart_1_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_system_burst_18_downstream_granted_uart_1_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_18_downstream_qualified_request_uart_1_s1 :  STD_LOGIC;
                signal internal_niosII_system_burst_18_downstream_requests_uart_1_s1 :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_arbiterlock :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_arbiterlock2 :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_continuerequest :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_saved_grant_uart_1_s1 :  STD_LOGIC;
                signal uart_1_s1_allgrants :  STD_LOGIC;
                signal uart_1_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal uart_1_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal uart_1_s1_any_continuerequest :  STD_LOGIC;
                signal uart_1_s1_arb_counter_enable :  STD_LOGIC;
                signal uart_1_s1_arb_share_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal uart_1_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal uart_1_s1_arb_share_set_values :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal uart_1_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal uart_1_s1_begins_xfer :  STD_LOGIC;
                signal uart_1_s1_end_xfer :  STD_LOGIC;
                signal uart_1_s1_firsttransfer :  STD_LOGIC;
                signal uart_1_s1_grant_vector :  STD_LOGIC;
                signal uart_1_s1_in_a_read_cycle :  STD_LOGIC;
                signal uart_1_s1_in_a_write_cycle :  STD_LOGIC;
                signal uart_1_s1_master_qreq_vector :  STD_LOGIC;
                signal uart_1_s1_non_bursting_master_requests :  STD_LOGIC;
                signal uart_1_s1_reg_firsttransfer :  STD_LOGIC;
                signal uart_1_s1_slavearbiterlockenable :  STD_LOGIC;
                signal uart_1_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal uart_1_s1_unreg_firsttransfer :  STD_LOGIC;
                signal uart_1_s1_waits_for_read :  STD_LOGIC;
                signal uart_1_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_uart_1_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT uart_1_s1_end_xfer;
    end if;

  end process;

  uart_1_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_system_burst_18_downstream_qualified_request_uart_1_s1);
  --assign uart_1_s1_readdata_from_sa = uart_1_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart_1_s1_readdata_from_sa <= uart_1_s1_readdata;
  internal_niosII_system_burst_18_downstream_requests_uart_1_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_system_burst_18_downstream_read OR niosII_system_burst_18_downstream_write)))))));
  --assign uart_1_s1_dataavailable_from_sa = uart_1_s1_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart_1_s1_dataavailable_from_sa <= uart_1_s1_dataavailable;
  --assign uart_1_s1_readyfordata_from_sa = uart_1_s1_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart_1_s1_readyfordata_from_sa <= uart_1_s1_readyfordata;
  --uart_1_s1_arb_share_counter set values, which is an e_mux
  uart_1_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_niosII_system_burst_18_downstream_granted_uart_1_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_18_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --uart_1_s1_non_bursting_master_requests mux, which is an e_mux
  uart_1_s1_non_bursting_master_requests <= std_logic'('0');
  --uart_1_s1_any_bursting_master_saved_grant mux, which is an e_mux
  uart_1_s1_any_bursting_master_saved_grant <= niosII_system_burst_18_downstream_saved_grant_uart_1_s1;
  --uart_1_s1_arb_share_counter_next_value assignment, which is an e_assign
  uart_1_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(uart_1_s1_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (uart_1_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(uart_1_s1_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000") & (uart_1_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 5);
  --uart_1_s1_allgrants all slave grants, which is an e_mux
  uart_1_s1_allgrants <= uart_1_s1_grant_vector;
  --uart_1_s1_end_xfer assignment, which is an e_assign
  uart_1_s1_end_xfer <= NOT ((uart_1_s1_waits_for_read OR uart_1_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_uart_1_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_uart_1_s1 <= uart_1_s1_end_xfer AND (((NOT uart_1_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --uart_1_s1_arb_share_counter arbitration counter enable, which is an e_assign
  uart_1_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_uart_1_s1 AND uart_1_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_uart_1_s1 AND NOT uart_1_s1_non_bursting_master_requests));
  --uart_1_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      uart_1_s1_arb_share_counter <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(uart_1_s1_arb_counter_enable) = '1' then 
        uart_1_s1_arb_share_counter <= uart_1_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --uart_1_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      uart_1_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((uart_1_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_uart_1_s1)) OR ((end_xfer_arb_share_counter_term_uart_1_s1 AND NOT uart_1_s1_non_bursting_master_requests)))) = '1' then 
        uart_1_s1_slavearbiterlockenable <= or_reduce(uart_1_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --niosII_system_burst_18/downstream uart_1/s1 arbiterlock, which is an e_assign
  niosII_system_burst_18_downstream_arbiterlock <= uart_1_s1_slavearbiterlockenable AND niosII_system_burst_18_downstream_continuerequest;
  --uart_1_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  uart_1_s1_slavearbiterlockenable2 <= or_reduce(uart_1_s1_arb_share_counter_next_value);
  --niosII_system_burst_18/downstream uart_1/s1 arbiterlock2, which is an e_assign
  niosII_system_burst_18_downstream_arbiterlock2 <= uart_1_s1_slavearbiterlockenable2 AND niosII_system_burst_18_downstream_continuerequest;
  --uart_1_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  uart_1_s1_any_continuerequest <= std_logic'('1');
  --niosII_system_burst_18_downstream_continuerequest continued request, which is an e_assign
  niosII_system_burst_18_downstream_continuerequest <= std_logic'('1');
  internal_niosII_system_burst_18_downstream_qualified_request_uart_1_s1 <= internal_niosII_system_burst_18_downstream_requests_uart_1_s1 AND NOT ((niosII_system_burst_18_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_18_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid niosII_system_burst_18_downstream_read_data_valid_uart_1_s1, which is an e_mux
  niosII_system_burst_18_downstream_read_data_valid_uart_1_s1 <= (internal_niosII_system_burst_18_downstream_granted_uart_1_s1 AND niosII_system_burst_18_downstream_read) AND NOT uart_1_s1_waits_for_read;
  --uart_1_s1_writedata mux, which is an e_mux
  uart_1_s1_writedata <= niosII_system_burst_18_downstream_writedata;
  --master is always granted when requested
  internal_niosII_system_burst_18_downstream_granted_uart_1_s1 <= internal_niosII_system_burst_18_downstream_qualified_request_uart_1_s1;
  --niosII_system_burst_18/downstream saved-grant uart_1/s1, which is an e_assign
  niosII_system_burst_18_downstream_saved_grant_uart_1_s1 <= internal_niosII_system_burst_18_downstream_requests_uart_1_s1;
  --allow new arb cycle for uart_1/s1, which is an e_assign
  uart_1_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  uart_1_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  uart_1_s1_master_qreq_vector <= std_logic'('1');
  uart_1_s1_begintransfer <= uart_1_s1_begins_xfer;
  --uart_1_s1_reset_n assignment, which is an e_assign
  uart_1_s1_reset_n <= reset_n;
  uart_1_s1_chipselect <= internal_niosII_system_burst_18_downstream_granted_uart_1_s1;
  --uart_1_s1_firsttransfer first transaction, which is an e_assign
  uart_1_s1_firsttransfer <= A_WE_StdLogic((std_logic'(uart_1_s1_begins_xfer) = '1'), uart_1_s1_unreg_firsttransfer, uart_1_s1_reg_firsttransfer);
  --uart_1_s1_unreg_firsttransfer first transaction, which is an e_assign
  uart_1_s1_unreg_firsttransfer <= NOT ((uart_1_s1_slavearbiterlockenable AND uart_1_s1_any_continuerequest));
  --uart_1_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      uart_1_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(uart_1_s1_begins_xfer) = '1' then 
        uart_1_s1_reg_firsttransfer <= uart_1_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --uart_1_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  uart_1_s1_beginbursttransfer_internal <= uart_1_s1_begins_xfer;
  --~uart_1_s1_read_n assignment, which is an e_mux
  uart_1_s1_read_n <= NOT ((internal_niosII_system_burst_18_downstream_granted_uart_1_s1 AND niosII_system_burst_18_downstream_read));
  --~uart_1_s1_write_n assignment, which is an e_mux
  uart_1_s1_write_n <= NOT ((internal_niosII_system_burst_18_downstream_granted_uart_1_s1 AND niosII_system_burst_18_downstream_write));
  --uart_1_s1_address mux, which is an e_mux
  uart_1_s1_address <= niosII_system_burst_18_downstream_nativeaddress (2 DOWNTO 0);
  --d1_uart_1_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_uart_1_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_uart_1_s1_end_xfer <= uart_1_s1_end_xfer;
    end if;

  end process;

  --uart_1_s1_waits_for_read in a cycle, which is an e_mux
  uart_1_s1_waits_for_read <= uart_1_s1_in_a_read_cycle AND uart_1_s1_begins_xfer;
  --uart_1_s1_in_a_read_cycle assignment, which is an e_assign
  uart_1_s1_in_a_read_cycle <= internal_niosII_system_burst_18_downstream_granted_uart_1_s1 AND niosII_system_burst_18_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= uart_1_s1_in_a_read_cycle;
  --uart_1_s1_waits_for_write in a cycle, which is an e_mux
  uart_1_s1_waits_for_write <= uart_1_s1_in_a_write_cycle AND uart_1_s1_begins_xfer;
  --uart_1_s1_in_a_write_cycle assignment, which is an e_assign
  uart_1_s1_in_a_write_cycle <= internal_niosII_system_burst_18_downstream_granted_uart_1_s1 AND niosII_system_burst_18_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= uart_1_s1_in_a_write_cycle;
  wait_for_uart_1_s1_counter <= std_logic'('0');
  --assign uart_1_s1_irq_from_sa = uart_1_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart_1_s1_irq_from_sa <= uart_1_s1_irq;
  --vhdl renameroo for output signals
  niosII_system_burst_18_downstream_granted_uart_1_s1 <= internal_niosII_system_burst_18_downstream_granted_uart_1_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_18_downstream_qualified_request_uart_1_s1 <= internal_niosII_system_burst_18_downstream_qualified_request_uart_1_s1;
  --vhdl renameroo for output signals
  niosII_system_burst_18_downstream_requests_uart_1_s1 <= internal_niosII_system_burst_18_downstream_requests_uart_1_s1;
--synthesis translate_off
    --uart_1/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --niosII_system_burst_18/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line220 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_18_downstream_requests_uart_1_s1 AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (niosII_system_burst_18_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line220, now);
          write(write_line220, string'(": "));
          write(write_line220, string'("niosII_system_burst_18/downstream drove 0 on its 'arbitrationshare' port while accessing slave uart_1/s1"));
          write(output, write_line220.all);
          deallocate (write_line220);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_system_burst_18/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line221 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_niosII_system_burst_18_downstream_requests_uart_1_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_system_burst_18_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line221, now);
          write(write_line221, string'(": "));
          write(write_line221, string'("niosII_system_burst_18/downstream drove 0 on its 'burstcount' port while accessing slave uart_1/s1"));
          write(output, write_line221.all);
          deallocate (write_line221);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_system_reset_clk_0_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity niosII_system_reset_clk_0_domain_synch_module;


architecture europa of niosII_system_reset_clk_0_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_system_reset_altpll_inst_c1_out_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity niosII_system_reset_altpll_inst_c1_out_domain_synch_module;


architecture europa of niosII_system_reset_altpll_inst_c1_out_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_system is 
        port (
              -- 1) global signals:
                 signal altpll_inst_c0_out : OUT STD_LOGIC;
                 signal altpll_inst_c1_out : OUT STD_LOGIC;
                 signal altpll_inst_c2_out : OUT STD_LOGIC;
                 signal clk_0 : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sram_IF_0_tsb_data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_altpll_inst
                 signal locked_from_the_altpll_inst : OUT STD_LOGIC;
                 signal phasedone_from_the_altpll_inst : OUT STD_LOGIC;

              -- the_dm9000a_inst
                 signal ENET_CMD_from_the_dm9000a_inst : OUT STD_LOGIC;
                 signal ENET_CS_N_from_the_dm9000a_inst : OUT STD_LOGIC;
                 signal ENET_DATA_to_and_from_the_dm9000a_inst : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal ENET_INT_to_the_dm9000a_inst : IN STD_LOGIC;
                 signal ENET_RD_N_from_the_dm9000a_inst : OUT STD_LOGIC;
                 signal ENET_RST_N_from_the_dm9000a_inst : OUT STD_LOGIC;
                 signal ENET_WR_N_from_the_dm9000a_inst : OUT STD_LOGIC;

              -- the_lcd_display
                 signal LCD_E_from_the_lcd_display : OUT STD_LOGIC;
                 signal LCD_RS_from_the_lcd_display : OUT STD_LOGIC;
                 signal LCD_RW_from_the_lcd_display : OUT STD_LOGIC;
                 signal LCD_data_to_and_from_the_lcd_display : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_led_pio
                 signal out_port_from_the_led_pio : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_sdram
                 signal zs_addr_from_the_sdram : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal zs_ba_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_cas_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_cke_from_the_sdram : OUT STD_LOGIC;
                 signal zs_cs_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_dq_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal zs_dqm_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_ras_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_we_n_from_the_sdram : OUT STD_LOGIC;

              -- the_seven_seg_pio
                 signal out_port_from_the_seven_seg_pio : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_sram_IF_0
                 signal coe_sram_address_from_the_sram_IF_0 : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal coe_sram_chipenable_n_from_the_sram_IF_0 : OUT STD_LOGIC;
                 signal coe_sram_lowerbyte_n_from_the_sram_IF_0 : OUT STD_LOGIC;
                 signal coe_sram_outputenable_n_from_the_sram_IF_0 : OUT STD_LOGIC;
                 signal coe_sram_upperbyte_n_from_the_sram_IF_0 : OUT STD_LOGIC;
                 signal coe_sram_writeenable_n_from_the_sram_IF_0 : OUT STD_LOGIC;

              -- the_switch
                 signal in_port_to_the_switch : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_tri_state_bridge_avalon_slave
                 signal address_to_the_ext_flash : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal data_to_and_from_the_ext_flash : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal read_n_to_the_ext_flash : OUT STD_LOGIC;
                 signal select_n_to_the_ext_flash : OUT STD_LOGIC;
                 signal write_n_to_the_ext_flash : OUT STD_LOGIC;

              -- the_uart_0
                 signal rxd_to_the_uart_0 : IN STD_LOGIC;
                 signal txd_from_the_uart_0 : OUT STD_LOGIC;

              -- the_uart_1
                 signal rxd_to_the_uart_1 : IN STD_LOGIC;
                 signal txd_from_the_uart_1 : OUT STD_LOGIC
              );
end entity niosII_system;


architecture europa of niosII_system is
component altpll_inst_pll_slave_arbitrator is 
           port (
                 -- inputs:
                    signal altpll_inst_pll_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_clock_0_out_read : IN STD_LOGIC;
                    signal niosII_system_clock_0_out_write : IN STD_LOGIC;
                    signal niosII_system_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal altpll_inst_pll_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal altpll_inst_pll_slave_read : OUT STD_LOGIC;
                    signal altpll_inst_pll_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal altpll_inst_pll_slave_reset : OUT STD_LOGIC;
                    signal altpll_inst_pll_slave_write : OUT STD_LOGIC;
                    signal altpll_inst_pll_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_altpll_inst_pll_slave_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_clock_0_out_granted_altpll_inst_pll_slave : OUT STD_LOGIC;
                    signal niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave : OUT STD_LOGIC;
                    signal niosII_system_clock_0_out_read_data_valid_altpll_inst_pll_slave : OUT STD_LOGIC;
                    signal niosII_system_clock_0_out_requests_altpll_inst_pll_slave : OUT STD_LOGIC
                 );
end component altpll_inst_pll_slave_arbitrator;

component altpll_inst is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal c0 : OUT STD_LOGIC;
                    signal c1 : OUT STD_LOGIC;
                    signal c2 : OUT STD_LOGIC;
                    signal locked : OUT STD_LOGIC;
                    signal phasedone : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component altpll_inst;

component cpu_jtag_debug_module_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_address_to_slave : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal niosII_system_burst_0_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_0_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_0_downstream_debugaccess : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_1_downstream_address_to_slave : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal niosII_system_burst_1_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_1_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_1_downstream_debugaccess : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal cpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_jtag_debug_module_reset_n : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_write : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_jtag_debug_module_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module : OUT STD_LOGIC
                 );
end component cpu_jtag_debug_module_arbitrator;

component cpu_data_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable_niosII_system_burst_11_upstream : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_byteenable_niosII_system_burst_13_upstream : IN STD_LOGIC;
                    signal cpu_data_master_byteenable_niosII_system_burst_20_upstream : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_granted_niosII_system_burst_11_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_13_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_14_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_15_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_16_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_17_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_18_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_1_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_20_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_21_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_3_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_4_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_5_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_6_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_7_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_8_upstream : IN STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_9_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_11_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_13_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_14_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_15_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_16_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_17_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_18_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_1_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_20_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_21_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_3_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_4_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_5_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_6_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_7_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_8_upstream : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_9_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_11_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_13_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_14_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_15_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_16_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_17_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_18_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_1_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_20_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_21_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_3_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_4_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_5_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_6_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_7_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_8_upstream : IN STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_9_upstream : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_niosII_system_burst_11_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_13_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_14_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_15_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_16_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_17_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_18_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_1_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_20_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_21_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_3_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_4_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_5_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_6_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_7_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_8_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_9_upstream_end_xfer : IN STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_irq_from_sa : IN STD_LOGIC;
                    signal high_res_timer_s1_irq_from_sa : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_11_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_11_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_13_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_13_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_14_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_14_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_15_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_15_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_16_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_16_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_17_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_17_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_18_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_18_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_1_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_1_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_20_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_20_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_21_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_21_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_3_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_3_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_4_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_4_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_5_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_5_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_6_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_6_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_7_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_7_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_8_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_8_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_9_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_9_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_timer_s1_irq_from_sa : IN STD_LOGIC;
                    signal uart_0_s1_irq_from_sa : IN STD_LOGIC;
                    signal uart_1_s1_irq_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal cpu_data_master_dbs_write_8 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal cpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_data_master_latency_counter : OUT STD_LOGIC;
                    signal cpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_data_master_readdatavalid : OUT STD_LOGIC;
                    signal cpu_data_master_waitrequest : OUT STD_LOGIC
                 );
end component cpu_data_master_arbitrator;

component cpu_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_instruction_master_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_instruction_master_granted_niosII_system_burst_0_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_granted_niosII_system_burst_10_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_granted_niosII_system_burst_12_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_granted_niosII_system_burst_19_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_granted_niosII_system_burst_2_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_requests_niosII_system_burst_0_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_requests_niosII_system_burst_10_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_requests_niosII_system_burst_12_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_requests_niosII_system_burst_19_upstream : IN STD_LOGIC;
                    signal cpu_instruction_master_requests_niosII_system_burst_2_upstream : IN STD_LOGIC;
                    signal d1_niosII_system_burst_0_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_10_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_12_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_19_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_system_burst_2_upstream_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_0_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_0_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_10_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_10_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_12_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_12_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_19_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_19_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_2_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_2_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : OUT STD_LOGIC;
                    signal cpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                    signal cpu_instruction_master_waitrequest : OUT STD_LOGIC
                 );
end component cpu_instruction_master_arbitrator;

component cpu is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d_irq : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdatavalid : IN STD_LOGIC;
                    signal d_waitrequest : IN STD_LOGIC;
                    signal i_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_readdatavalid : IN STD_LOGIC;
                    signal i_waitrequest : IN STD_LOGIC;
                    signal jtag_debug_module_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal jtag_debug_module_begintransfer : IN STD_LOGIC;
                    signal jtag_debug_module_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal jtag_debug_module_debugaccess : IN STD_LOGIC;
                    signal jtag_debug_module_select : IN STD_LOGIC;
                    signal jtag_debug_module_write : IN STD_LOGIC;
                    signal jtag_debug_module_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal d_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_read : OUT STD_LOGIC;
                    signal d_write : OUT STD_LOGIC;
                    signal d_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal i_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal i_read : OUT STD_LOGIC;
                    signal jtag_debug_module_debugaccess_to_roms : OUT STD_LOGIC;
                    signal jtag_debug_module_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_debug_module_resetrequest : OUT STD_LOGIC
                 );
end component cpu;

component dm9000a_inst_avalon_slave_0_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_irq : IN STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_16_downstream_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_16_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_16_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_16_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_dm9000a_inst_avalon_slave_0_end_xfer : OUT STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_address : OUT STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_chipselect_n : OUT STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_irq_from_sa : OUT STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_read_n : OUT STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal dm9000a_inst_avalon_slave_0_reset_n : OUT STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_write_n : OUT STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 : OUT STD_LOGIC;
                    signal niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 : OUT STD_LOGIC;
                    signal niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0 : OUT STD_LOGIC;
                    signal niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 : OUT STD_LOGIC
                 );
end component dm9000a_inst_avalon_slave_0_arbitrator;

component dm9000a_inst is 
           port (
                 -- inputs:
                    signal ENET_INT : IN STD_LOGIC;
                    signal iCMD : IN STD_LOGIC;
                    signal iCS_N : IN STD_LOGIC;
                    signal iDATA : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal iRD_N : IN STD_LOGIC;
                    signal iRST_N : IN STD_LOGIC;
                    signal iWR_N : IN STD_LOGIC;

                 -- outputs:
                    signal ENET_CMD : OUT STD_LOGIC;
                    signal ENET_CS_N : OUT STD_LOGIC;
                    signal ENET_DATA : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal ENET_RD_N : OUT STD_LOGIC;
                    signal ENET_RST_N : OUT STD_LOGIC;
                    signal ENET_WR_N : OUT STD_LOGIC;
                    signal oDATA : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal oINT : OUT STD_LOGIC
                 );
end component dm9000a_inst;

component high_res_timer_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal high_res_timer_s1_irq : IN STD_LOGIC;
                    signal high_res_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_15_downstream_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_15_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_15_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_15_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_high_res_timer_s1_end_xfer : OUT STD_LOGIC;
                    signal high_res_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal high_res_timer_s1_chipselect : OUT STD_LOGIC;
                    signal high_res_timer_s1_irq_from_sa : OUT STD_LOGIC;
                    signal high_res_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal high_res_timer_s1_reset_n : OUT STD_LOGIC;
                    signal high_res_timer_s1_write_n : OUT STD_LOGIC;
                    signal high_res_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_15_downstream_granted_high_res_timer_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_15_downstream_requests_high_res_timer_s1 : OUT STD_LOGIC
                 );
end component high_res_timer_s1_arbitrator;

component high_res_timer is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component high_res_timer;

component jtag_uart_avalon_jtag_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_6_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_6_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_6_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC
                 );
end component jtag_uart_avalon_jtag_slave_arbitrator;

component jtag_uart is 
           port (
                 -- inputs:
                    signal av_address : IN STD_LOGIC;
                    signal av_chipselect : IN STD_LOGIC;
                    signal av_read_n : IN STD_LOGIC;
                    signal av_write_n : IN STD_LOGIC;
                    signal av_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_irq : OUT STD_LOGIC;
                    signal av_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_waitrequest : OUT STD_LOGIC;
                    signal dataavailable : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component jtag_uart;

component lcd_display_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_display_control_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_7_downstream_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_7_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal niosII_system_burst_7_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_byteenable : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_7_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_lcd_display_control_slave_end_xfer : OUT STD_LOGIC;
                    signal lcd_display_control_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_display_control_slave_begintransfer : OUT STD_LOGIC;
                    signal lcd_display_control_slave_read : OUT STD_LOGIC;
                    signal lcd_display_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal lcd_display_control_slave_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal lcd_display_control_slave_write : OUT STD_LOGIC;
                    signal lcd_display_control_slave_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_7_downstream_granted_lcd_display_control_slave : OUT STD_LOGIC;
                    signal niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave : OUT STD_LOGIC;
                    signal niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave : OUT STD_LOGIC;
                    signal niosII_system_burst_7_downstream_requests_lcd_display_control_slave : OUT STD_LOGIC
                 );
end component lcd_display_control_slave_arbitrator;

component lcd_display is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal begintransfer : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal LCD_E : OUT STD_LOGIC;
                    signal LCD_RS : OUT STD_LOGIC;
                    signal LCD_RW : OUT STD_LOGIC;
                    signal LCD_data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component lcd_display;

component led_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal led_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_8_downstream_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_8_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal niosII_system_burst_8_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_byteenable : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_8_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_led_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal led_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal led_pio_s1_chipselect : OUT STD_LOGIC;
                    signal led_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal led_pio_s1_reset_n : OUT STD_LOGIC;
                    signal led_pio_s1_write_n : OUT STD_LOGIC;
                    signal led_pio_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_8_downstream_granted_led_pio_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_8_downstream_qualified_request_led_pio_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_8_downstream_read_data_valid_led_pio_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_8_downstream_requests_led_pio_s1 : OUT STD_LOGIC
                 );
end component led_pio_s1_arbitrator;

component led_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component led_pio;

component memory_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_2_downstream_address_to_slave : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal niosII_system_burst_2_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_2_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_2_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_3_downstream_address_to_slave : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal niosII_system_burst_3_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_3_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_3_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_memory_s1_end_xfer : OUT STD_LOGIC;
                    signal memory_s1_address : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal memory_s1_chipselect : OUT STD_LOGIC;
                    signal memory_s1_clken : OUT STD_LOGIC;
                    signal memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal memory_s1_reset : OUT STD_LOGIC;
                    signal memory_s1_write : OUT STD_LOGIC;
                    signal memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_2_downstream_granted_memory_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_2_downstream_qualified_request_memory_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_2_downstream_read_data_valid_memory_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_2_downstream_requests_memory_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_3_downstream_granted_memory_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_3_downstream_qualified_request_memory_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_3_downstream_read_data_valid_memory_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_3_downstream_requests_memory_s1 : OUT STD_LOGIC
                 );
end component memory_s1_arbitrator;

component memory is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clken : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component memory;

component niosII_system_burst_0_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : IN STD_LOGIC;
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : IN STD_LOGIC;
                    signal niosII_system_burst_0_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_0_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_0_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_instruction_master_granted_niosII_system_burst_0_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_instruction_master_requests_niosII_system_burst_0_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_0_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_0_upstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal niosII_system_burst_0_upstream_byteaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal niosII_system_burst_0_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_0_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_0_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_0_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_0_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_0_upstream_write : OUT STD_LOGIC
                 );
end component niosII_system_burst_0_upstream_arbitrator;

component niosII_system_burst_0_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal niosII_system_burst_0_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_0_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal niosII_system_burst_0_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_0_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_0_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_0_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_0_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_0_downstream_arbitrator;

component niosII_system_burst_0 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_0;

component niosII_system_burst_1_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_1_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_1_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_1_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_1_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_1_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_1_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_1_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_1_upstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal niosII_system_burst_1_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_1_upstream_byteaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal niosII_system_burst_1_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_1_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_1_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_1_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_1_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_1_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_1_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component niosII_system_burst_1_upstream_arbitrator;

component niosII_system_burst_1_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal niosII_system_burst_1_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_1_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal niosII_system_burst_1_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_1_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_1_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_1_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_1_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_1_downstream_arbitrator;

component niosII_system_burst_1 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_1;

component niosII_system_burst_10_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : IN STD_LOGIC;
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : IN STD_LOGIC;
                    signal niosII_system_burst_10_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_10_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_10_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_instruction_master_granted_niosII_system_burst_10_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_instruction_master_requests_niosII_system_burst_10_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_10_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_10_upstream_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal niosII_system_burst_10_upstream_byteaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal niosII_system_burst_10_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_10_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_10_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_10_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_10_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_10_upstream_write : OUT STD_LOGIC
                 );
end component niosII_system_burst_10_upstream_arbitrator;

component niosII_system_burst_10_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal niosII_system_burst_10_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_10_downstream_granted_sdram_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_requests_sdram_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_10_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal niosII_system_burst_10_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_10_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_10_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_10_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_10_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_10_downstream_arbitrator;

component niosII_system_burst_10 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_10;

component niosII_system_burst_11_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal niosII_system_burst_11_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_11_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_11_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_byteenable_niosII_system_burst_11_upstream : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_granted_niosII_system_burst_11_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_11_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_11_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_11_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_11_upstream_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal niosII_system_burst_11_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_11_upstream_byteaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal niosII_system_burst_11_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_11_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_11_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_11_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_11_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_11_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_11_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component niosII_system_burst_11_upstream_arbitrator;

component niosII_system_burst_11_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal niosII_system_burst_11_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_11_downstream_granted_sdram_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_requests_sdram_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_11_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal niosII_system_burst_11_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_11_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_11_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_11_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_11_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_11_downstream_arbitrator;

component niosII_system_burst_11 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_11;

component niosII_system_burst_12_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : IN STD_LOGIC;
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : IN STD_LOGIC;
                    signal niosII_system_burst_12_upstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_12_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_12_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_instruction_master_granted_niosII_system_burst_12_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_instruction_master_requests_niosII_system_burst_12_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_12_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_12_upstream_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal niosII_system_burst_12_upstream_byteaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal niosII_system_burst_12_upstream_byteenable : OUT STD_LOGIC;
                    signal niosII_system_burst_12_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_12_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_12_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_12_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_12_upstream_write : OUT STD_LOGIC
                 );
end component niosII_system_burst_12_upstream_arbitrator;

component niosII_system_burst_12_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_tri_state_bridge_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal ext_flash_s1_wait_counter_eq_0 : IN STD_LOGIC;
                    signal incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_12_downstream_address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal niosII_system_burst_12_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_byteenable : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_granted_ext_flash_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_requests_ext_flash_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_12_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal niosII_system_burst_12_downstream_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_12_downstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_12_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_12_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_12_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_12_downstream_arbitrator;

component niosII_system_burst_12 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC;
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC;
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_12;

component niosII_system_burst_13_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal niosII_system_burst_13_upstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_13_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_13_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_byteenable_niosII_system_burst_13_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_granted_niosII_system_burst_13_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_13_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_13_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_13_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_13_upstream_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal niosII_system_burst_13_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_13_upstream_byteaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal niosII_system_burst_13_upstream_byteenable : OUT STD_LOGIC;
                    signal niosII_system_burst_13_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_13_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_13_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_13_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_13_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_13_upstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component niosII_system_burst_13_upstream_arbitrator;

component niosII_system_burst_13_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_tri_state_bridge_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal ext_flash_s1_wait_counter_eq_0 : IN STD_LOGIC;
                    signal incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_13_downstream_address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal niosII_system_burst_13_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_byteenable : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_granted_ext_flash_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_requests_ext_flash_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_13_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal niosII_system_burst_13_downstream_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_13_downstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_13_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_13_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_13_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_13_downstream_arbitrator;

component niosII_system_burst_13 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC;
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC;
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_13;

component niosII_system_burst_14_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_14_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_14_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_14_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_14_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_14_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_14_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_14_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_14_upstream_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_14_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_14_upstream_byteaddress : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_14_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_14_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_14_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_14_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_14_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_14_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_14_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component niosII_system_burst_14_upstream_arbitrator;

component niosII_system_burst_14_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_seven_seg_pio_s1_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_14_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal seven_seg_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal niosII_system_burst_14_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_14_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_14_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_14_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_14_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_14_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_14_downstream_arbitrator;

component niosII_system_burst_14 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_14;

component niosII_system_burst_15_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_15_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_15_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_15_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_15_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_15_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_15_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_15_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_15_upstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_15_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_15_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_15_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_15_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_15_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_15_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_15_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_15_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_15_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component niosII_system_burst_15_upstream_arbitrator;

component niosII_system_burst_15_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_high_res_timer_s1_end_xfer : IN STD_LOGIC;
                    signal high_res_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_15_downstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_15_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_15_downstream_granted_high_res_timer_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_requests_high_res_timer_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_15_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_15_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_15_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_15_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_15_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_15_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_15_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_15_downstream_arbitrator;

component niosII_system_burst_15 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_15;

component niosII_system_burst_16_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_16_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_16_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_16_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_16_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_16_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_16_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_16_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_16_upstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_16_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_16_upstream_byteaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_16_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_16_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_16_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_16_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_16_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_16_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_16_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component niosII_system_burst_16_upstream_arbitrator;

component niosII_system_burst_16_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_dm9000a_inst_avalon_slave_0_end_xfer : IN STD_LOGIC;
                    signal dm9000a_inst_avalon_slave_0_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_16_downstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_16_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0 : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_16_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_16_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_16_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_16_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_16_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_16_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_16_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_16_downstream_arbitrator;

component niosII_system_burst_16 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_16;

component niosII_system_burst_17_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_17_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_17_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_17_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_17_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_17_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_17_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_17_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_17_upstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_17_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_17_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_17_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_17_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_17_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_17_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_17_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_17_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_17_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component niosII_system_burst_17_upstream_arbitrator;

component niosII_system_burst_17_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_uart_0_s1_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_17_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_17_downstream_granted_uart_0_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_qualified_request_uart_0_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_read_data_valid_uart_0_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_requests_uart_0_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal uart_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal niosII_system_burst_17_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_17_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_17_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_17_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_17_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_17_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_17_downstream_arbitrator;

component niosII_system_burst_17 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_17;

component niosII_system_burst_18_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_18_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_18_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_18_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_18_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_18_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_18_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_18_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_18_upstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_18_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_18_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_18_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_18_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_18_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_18_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_18_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_18_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_18_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component niosII_system_burst_18_upstream_arbitrator;

component niosII_system_burst_18_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_uart_1_s1_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_18_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_18_downstream_granted_uart_1_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_qualified_request_uart_1_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_read_data_valid_uart_1_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_requests_uart_1_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal uart_1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal niosII_system_burst_18_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_18_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_18_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_18_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_18_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_18_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_18_downstream_arbitrator;

component niosII_system_burst_18 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_18;

component niosII_system_burst_19_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : IN STD_LOGIC;
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : IN STD_LOGIC;
                    signal niosII_system_burst_19_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_19_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_19_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_instruction_master_granted_niosII_system_burst_19_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_instruction_master_requests_niosII_system_burst_19_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_19_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_19_upstream_address : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal niosII_system_burst_19_upstream_byteaddress : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
                    signal niosII_system_burst_19_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_19_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_19_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_19_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_19_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_19_upstream_write : OUT STD_LOGIC
                 );
end component niosII_system_burst_19_upstream_arbitrator;

component niosII_system_burst_19_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_tsb_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal incoming_sram_IF_0_tsb_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_address : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_granted_sram_IF_0_tsb : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_requests_sram_IF_0_tsb : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_19_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_19_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_19_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_19_downstream_arbitrator;

component niosII_system_burst_19 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (19 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_19;

component niosII_system_burst_2_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : IN STD_LOGIC;
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register : IN STD_LOGIC;
                    signal niosII_system_burst_2_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_2_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_2_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_instruction_master_granted_niosII_system_burst_2_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_instruction_master_requests_niosII_system_burst_2_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_2_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_2_upstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal niosII_system_burst_2_upstream_byteaddress : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_2_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_2_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_2_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_2_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_2_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_2_upstream_write : OUT STD_LOGIC
                 );
end component niosII_system_burst_2_upstream_arbitrator;

component niosII_system_burst_2_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_memory_s1_end_xfer : IN STD_LOGIC;
                    signal memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_2_downstream_address : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal niosII_system_burst_2_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_2_downstream_granted_memory_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_qualified_request_memory_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_read_data_valid_memory_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_requests_memory_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_2_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal niosII_system_burst_2_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_2_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_2_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_2_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_2_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_2_downstream_arbitrator;

component niosII_system_burst_2 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_2;

component niosII_system_burst_20_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal niosII_system_burst_20_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_20_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_20_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_byteenable_niosII_system_burst_20_upstream : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_granted_niosII_system_burst_20_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_20_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_20_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_20_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_20_upstream_address : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal niosII_system_burst_20_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_20_upstream_byteaddress : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
                    signal niosII_system_burst_20_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_20_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_20_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_20_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_20_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_20_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_20_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component niosII_system_burst_20_upstream_arbitrator;

component niosII_system_burst_20_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_tsb_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal incoming_sram_IF_0_tsb_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_address : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_20_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_granted_sram_IF_0_tsb : IN STD_LOGIC;
                    signal niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb : IN STD_LOGIC;
                    signal niosII_system_burst_20_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb : IN STD_LOGIC;
                    signal niosII_system_burst_20_downstream_requests_sram_IF_0_tsb : IN STD_LOGIC;
                    signal niosII_system_burst_20_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_20_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_20_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_20_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_20_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_20_downstream_arbitrator;

component niosII_system_burst_20 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (19 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_20;

component niosII_system_burst_21_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_21_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_21_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_21_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_21_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_21_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_21_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_21_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_21_upstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_21_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_21_upstream_byteaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal niosII_system_burst_21_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_21_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_21_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_21_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_21_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_21_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_21_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component niosII_system_burst_21_upstream_arbitrator;

component niosII_system_burst_21_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_niosII_system_clock_0_in_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_21_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_21_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_21_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_21_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_21_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_21_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_21_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_21_downstream_arbitrator;

component niosII_system_burst_21 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_21;

component niosII_system_burst_3_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_3_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_3_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_3_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_3_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_3_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_3_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_3_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_3_upstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal niosII_system_burst_3_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_3_upstream_byteaddress : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_3_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_3_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_3_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_3_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_3_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_3_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_3_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component niosII_system_burst_3_upstream_arbitrator;

component niosII_system_burst_3_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_memory_s1_end_xfer : IN STD_LOGIC;
                    signal memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_3_downstream_address : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal niosII_system_burst_3_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_3_downstream_granted_memory_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_qualified_request_memory_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_read_data_valid_memory_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_requests_memory_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_3_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal niosII_system_burst_3_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_3_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_3_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_3_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_3_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_3_downstream_arbitrator;

component niosII_system_burst_3 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_3;

component niosII_system_burst_4_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_4_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_4_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_4_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_4_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_4_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_4_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_4_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_4_upstream_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_4_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_4_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_4_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_4_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_4_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_4_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_4_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_4_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_4_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component niosII_system_burst_4_upstream_arbitrator;

component niosII_system_burst_4_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_4_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_4_downstream_granted_sysid_control_slave : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_qualified_request_sysid_control_slave : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_requests_sysid_control_slave : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal niosII_system_burst_4_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_4_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_4_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_4_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_4_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_4_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_4_downstream_arbitrator;

component niosII_system_burst_4 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_4;

component niosII_system_burst_5_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_5_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_5_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_5_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_5_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_5_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_5_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_5_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_5_upstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_5_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_5_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_5_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_5_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_5_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_5_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_5_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_5_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_5_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component niosII_system_burst_5_upstream_arbitrator;

component niosII_system_burst_5_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sys_clk_timer_s1_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_5_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal niosII_system_burst_5_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_5_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_5_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_5_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_5_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_5_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_5_downstream_arbitrator;

component niosII_system_burst_5 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_5;

component niosII_system_burst_6_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_6_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_6_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_6_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_6_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_6_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_6_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_6_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_6_upstream_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_6_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_6_upstream_byteaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_6_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_6_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_6_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_6_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_6_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_6_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_6_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component niosII_system_burst_6_upstream_arbitrator;

component niosII_system_burst_6_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_6_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_6_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_6_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_6_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_6_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_6_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_6_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_6_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_6_downstream_arbitrator;

component niosII_system_burst_6 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_6;

component niosII_system_burst_7_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_7_upstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_7_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_7_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_7_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_7_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_7_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_7_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_7_upstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_7_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_7_upstream_byteaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_7_upstream_byteenable : OUT STD_LOGIC;
                    signal niosII_system_burst_7_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_7_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_7_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_7_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_7_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_7_upstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component niosII_system_burst_7_upstream_arbitrator;

component niosII_system_burst_7_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_lcd_display_control_slave_end_xfer : IN STD_LOGIC;
                    signal lcd_display_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal lcd_display_control_slave_wait_counter_eq_0 : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_7_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_byteenable : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_granted_lcd_display_control_slave : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_requests_lcd_display_control_slave : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_7_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_7_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_7_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_7_downstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_7_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_7_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_7_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_7_downstream_arbitrator;

component niosII_system_burst_7 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC;
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC;
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_7;

component niosII_system_burst_8_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_8_upstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_8_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_8_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_8_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_8_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_8_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_8_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_8_upstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_8_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_8_upstream_byteaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_8_upstream_byteenable : OUT STD_LOGIC;
                    signal niosII_system_burst_8_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_8_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_8_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_8_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_8_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_8_upstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component niosII_system_burst_8_upstream_arbitrator;

component niosII_system_burst_8_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_led_pio_s1_end_xfer : IN STD_LOGIC;
                    signal led_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_8_downstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_8_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_byteenable : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_granted_led_pio_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_qualified_request_led_pio_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_read_data_valid_led_pio_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_requests_led_pio_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_8_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_burst_8_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_8_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_8_downstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_8_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_8_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_8_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_8_downstream_arbitrator;

component niosII_system_burst_8 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC;
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC;
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_8;

component niosII_system_burst_9_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_burst_9_upstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_9_upstream_readdatavalid : IN STD_LOGIC;
                    signal niosII_system_burst_9_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_niosII_system_burst_9_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_niosII_system_burst_9_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_niosII_system_burst_9_upstream : OUT STD_LOGIC;
                    signal d1_niosII_system_burst_9_upstream_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_9_upstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_9_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_9_upstream_byteaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_9_upstream_byteenable : OUT STD_LOGIC;
                    signal niosII_system_burst_9_upstream_debugaccess : OUT STD_LOGIC;
                    signal niosII_system_burst_9_upstream_read : OUT STD_LOGIC;
                    signal niosII_system_burst_9_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_9_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_burst_9_upstream_write : OUT STD_LOGIC;
                    signal niosII_system_burst_9_upstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component niosII_system_burst_9_upstream_arbitrator;

component niosII_system_burst_9_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_switch_s1_end_xfer : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_9_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_byteenable : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_granted_switch_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_qualified_request_switch_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_read_data_valid_switch_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_requests_switch_s1 : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal switch_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal niosII_system_burst_9_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_9_downstream_latency_counter : OUT STD_LOGIC;
                    signal niosII_system_burst_9_downstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_9_downstream_readdatavalid : OUT STD_LOGIC;
                    signal niosII_system_burst_9_downstream_reset_n : OUT STD_LOGIC;
                    signal niosII_system_burst_9_downstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_9_downstream_arbitrator;

component niosII_system_burst_9 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC;
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC;
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_burst_9;

component niosII_system_clock_0_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_21_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_21_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_21_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_21_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_21_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_clock_0_in_endofpacket : IN STD_LOGIC;
                    signal niosII_system_clock_0_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_clock_0_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_niosII_system_clock_0_in_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in : OUT STD_LOGIC;
                    signal niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in : OUT STD_LOGIC;
                    signal niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in : OUT STD_LOGIC;
                    signal niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in : OUT STD_LOGIC;
                    signal niosII_system_clock_0_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal niosII_system_clock_0_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_clock_0_in_read : OUT STD_LOGIC;
                    signal niosII_system_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_clock_0_in_reset_n : OUT STD_LOGIC;
                    signal niosII_system_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_system_clock_0_in_write : OUT STD_LOGIC;
                    signal niosII_system_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component niosII_system_clock_0_in_arbitrator;

component niosII_system_clock_0_out_arbitrator is 
           port (
                 -- inputs:
                    signal altpll_inst_pll_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_altpll_inst_pll_slave_end_xfer : IN STD_LOGIC;
                    signal niosII_system_clock_0_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_clock_0_out_granted_altpll_inst_pll_slave : IN STD_LOGIC;
                    signal niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave : IN STD_LOGIC;
                    signal niosII_system_clock_0_out_read : IN STD_LOGIC;
                    signal niosII_system_clock_0_out_read_data_valid_altpll_inst_pll_slave : IN STD_LOGIC;
                    signal niosII_system_clock_0_out_requests_altpll_inst_pll_slave : IN STD_LOGIC;
                    signal niosII_system_clock_0_out_write : IN STD_LOGIC;
                    signal niosII_system_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_system_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_system_clock_0_out_reset_n : OUT STD_LOGIC;
                    signal niosII_system_clock_0_out_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_clock_0_out_arbitrator;

component niosII_system_clock_0 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component niosII_system_clock_0;

component sdram_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_address_to_slave : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal niosII_system_burst_10_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_10_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_10_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_10_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_11_downstream_address_to_slave : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal niosII_system_burst_11_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_11_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_11_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_11_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_readdatavalid : IN STD_LOGIC;
                    signal sdram_s1_waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal d1_sdram_s1_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_10_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_10_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_10_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_10_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal niosII_system_burst_10_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_11_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_11_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_11_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_11_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal niosII_system_burst_11_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                    signal sdram_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal sdram_s1_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sdram_s1_chipselect : OUT STD_LOGIC;
                    signal sdram_s1_read_n : OUT STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_reset_n : OUT STD_LOGIC;
                    signal sdram_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal sdram_s1_write_n : OUT STD_LOGIC;
                    signal sdram_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sdram_s1_arbitrator;

component sdram is 
           port (
                 -- inputs:
                    signal az_addr : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal az_be_n : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal az_cs : IN STD_LOGIC;
                    signal az_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal az_rd_n : IN STD_LOGIC;
                    signal az_wr_n : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal za_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal za_valid : OUT STD_LOGIC;
                    signal za_waitrequest : OUT STD_LOGIC;
                    signal zs_addr : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n : OUT STD_LOGIC;
                    signal zs_cke : OUT STD_LOGIC;
                    signal zs_cs_n : OUT STD_LOGIC;
                    signal zs_dq : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal zs_dqm : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n : OUT STD_LOGIC;
                    signal zs_we_n : OUT STD_LOGIC
                 );
end component sdram;

component seven_seg_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_14_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_14_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_14_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_14_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal seven_seg_pio_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal d1_seven_seg_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 : OUT STD_LOGIC;
                    signal seven_seg_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal seven_seg_pio_s1_chipselect : OUT STD_LOGIC;
                    signal seven_seg_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal seven_seg_pio_s1_reset_n : OUT STD_LOGIC;
                    signal seven_seg_pio_s1_write_n : OUT STD_LOGIC;
                    signal seven_seg_pio_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component seven_seg_pio_s1_arbitrator;

component seven_seg_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component seven_seg_pio;

component sram_IF_0 is 
           port (
                 -- inputs:
                    signal ats_tsb_address : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal ats_tsb_byteenable_n : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ats_tsb_chipselect_n : IN STD_LOGIC;
                    signal ats_tsb_outputenable_n : IN STD_LOGIC;
                    signal ats_tsb_write_n : IN STD_LOGIC;

                 -- outputs:
                    signal ats_tsb_data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal coe_sram_address : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal coe_sram_chipenable_n : OUT STD_LOGIC;
                    signal coe_sram_lowerbyte_n : OUT STD_LOGIC;
                    signal coe_sram_outputenable_n : OUT STD_LOGIC;
                    signal coe_sram_upperbyte_n : OUT STD_LOGIC;
                    signal coe_sram_writeenable_n : OUT STD_LOGIC
                 );
end component sram_IF_0;

component switch_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_9_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal niosII_system_burst_9_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_9_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_9_downstream_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal switch_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal d1_switch_s1_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_9_downstream_granted_switch_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_9_downstream_qualified_request_switch_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_9_downstream_read_data_valid_switch_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_9_downstream_requests_switch_s1 : OUT STD_LOGIC;
                    signal switch_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal switch_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal switch_s1_reset_n : OUT STD_LOGIC
                 );
end component switch_s1_arbitrator;

component switch is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component switch;

component sys_clk_timer_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_5_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_5_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_5_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_timer_s1_irq : IN STD_LOGIC;
                    signal sys_clk_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal d1_sys_clk_timer_s1_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal sys_clk_timer_s1_chipselect : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_irq_from_sa : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sys_clk_timer_s1_reset_n : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_write_n : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sys_clk_timer_s1_arbitrator;

component sys_clk_timer is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sys_clk_timer;

component sysid_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_4_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_4_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_system_burst_4_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_4_downstream_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_4_downstream_granted_sysid_control_slave : OUT STD_LOGIC;
                    signal niosII_system_burst_4_downstream_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                    signal niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                    signal niosII_system_burst_4_downstream_requests_sysid_control_slave : OUT STD_LOGIC;
                    signal sysid_control_slave_address : OUT STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sysid_control_slave_reset_n : OUT STD_LOGIC
                 );
end component sysid_control_slave_arbitrator;

component sysid is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC;
                    signal clock : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sysid;

component tri_state_bridge_avalon_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_address_to_slave : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal niosII_system_burst_12_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal niosII_system_burst_12_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_byteenable : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_12_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_12_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_13_downstream_address_to_slave : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal niosII_system_burst_13_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal niosII_system_burst_13_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_byteenable : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_13_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_13_downstream_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal address_to_the_ext_flash : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal d1_tri_state_bridge_avalon_slave_end_xfer : OUT STD_LOGIC;
                    signal data_to_and_from_the_ext_flash : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal ext_flash_s1_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_system_burst_12_downstream_granted_ext_flash_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_12_downstream_requests_ext_flash_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_13_downstream_granted_ext_flash_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_13_downstream_requests_ext_flash_s1 : OUT STD_LOGIC;
                    signal read_n_to_the_ext_flash : OUT STD_LOGIC;
                    signal select_n_to_the_ext_flash : OUT STD_LOGIC;
                    signal write_n_to_the_ext_flash : OUT STD_LOGIC
                 );
end component tri_state_bridge_avalon_slave_arbitrator;

component tri_state_bridge is 
end component tri_state_bridge;

component tri_state_bridge_bridge_arbitrator is 
end component tri_state_bridge_bridge_arbitrator;

component tsb_avalon_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_address_to_slave : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_19_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_address_to_slave : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_20_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_system_burst_20_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_20_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_20_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_tsb_avalon_slave_end_xfer : OUT STD_LOGIC;
                    signal incoming_sram_IF_0_tsb_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_system_burst_19_downstream_granted_sram_IF_0_tsb : OUT STD_LOGIC;
                    signal niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb : OUT STD_LOGIC;
                    signal niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb : OUT STD_LOGIC;
                    signal niosII_system_burst_19_downstream_requests_sram_IF_0_tsb : OUT STD_LOGIC;
                    signal niosII_system_burst_20_downstream_granted_sram_IF_0_tsb : OUT STD_LOGIC;
                    signal niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb : OUT STD_LOGIC;
                    signal niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb : OUT STD_LOGIC;
                    signal niosII_system_burst_20_downstream_requests_sram_IF_0_tsb : OUT STD_LOGIC;
                    signal sram_IF_0_tsb_address : OUT STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal sram_IF_0_tsb_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sram_IF_0_tsb_chipselect_n : OUT STD_LOGIC;
                    signal sram_IF_0_tsb_data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sram_IF_0_tsb_outputenable_n : OUT STD_LOGIC;
                    signal sram_IF_0_tsb_write_n : OUT STD_LOGIC
                 );
end component tsb_avalon_slave_arbitrator;

component tsb is 
end component tsb;

component tsb_bridge_arbitrator is 
end component tsb_bridge_arbitrator;

component uart_0_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_17_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_17_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_17_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_17_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal uart_0_s1_dataavailable : IN STD_LOGIC;
                    signal uart_0_s1_irq : IN STD_LOGIC;
                    signal uart_0_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal uart_0_s1_readyfordata : IN STD_LOGIC;

                 -- outputs:
                    signal d1_uart_0_s1_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_17_downstream_granted_uart_0_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_17_downstream_qualified_request_uart_0_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_17_downstream_read_data_valid_uart_0_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_17_downstream_requests_uart_0_s1 : OUT STD_LOGIC;
                    signal uart_0_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal uart_0_s1_begintransfer : OUT STD_LOGIC;
                    signal uart_0_s1_chipselect : OUT STD_LOGIC;
                    signal uart_0_s1_dataavailable_from_sa : OUT STD_LOGIC;
                    signal uart_0_s1_irq_from_sa : OUT STD_LOGIC;
                    signal uart_0_s1_read_n : OUT STD_LOGIC;
                    signal uart_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal uart_0_s1_readyfordata_from_sa : OUT STD_LOGIC;
                    signal uart_0_s1_reset_n : OUT STD_LOGIC;
                    signal uart_0_s1_write_n : OUT STD_LOGIC;
                    signal uart_0_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component uart_0_s1_arbitrator;

component uart_0 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal begintransfer : IN STD_LOGIC;
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal rxd : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal dataavailable : OUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readyfordata : OUT STD_LOGIC;
                    signal txd : OUT STD_LOGIC
                 );
end component uart_0;

component uart_1_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_18_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal niosII_system_burst_18_downstream_burstcount : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_latency_counter : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_nativeaddress : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_system_burst_18_downstream_read : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_write : IN STD_LOGIC;
                    signal niosII_system_burst_18_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal uart_1_s1_dataavailable : IN STD_LOGIC;
                    signal uart_1_s1_irq : IN STD_LOGIC;
                    signal uart_1_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal uart_1_s1_readyfordata : IN STD_LOGIC;

                 -- outputs:
                    signal d1_uart_1_s1_end_xfer : OUT STD_LOGIC;
                    signal niosII_system_burst_18_downstream_granted_uart_1_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_18_downstream_qualified_request_uart_1_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_18_downstream_read_data_valid_uart_1_s1 : OUT STD_LOGIC;
                    signal niosII_system_burst_18_downstream_requests_uart_1_s1 : OUT STD_LOGIC;
                    signal uart_1_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal uart_1_s1_begintransfer : OUT STD_LOGIC;
                    signal uart_1_s1_chipselect : OUT STD_LOGIC;
                    signal uart_1_s1_dataavailable_from_sa : OUT STD_LOGIC;
                    signal uart_1_s1_irq_from_sa : OUT STD_LOGIC;
                    signal uart_1_s1_read_n : OUT STD_LOGIC;
                    signal uart_1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal uart_1_s1_readyfordata_from_sa : OUT STD_LOGIC;
                    signal uart_1_s1_reset_n : OUT STD_LOGIC;
                    signal uart_1_s1_write_n : OUT STD_LOGIC;
                    signal uart_1_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component uart_1_s1_arbitrator;

component uart_1 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal begintransfer : IN STD_LOGIC;
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal rxd : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal dataavailable : OUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readyfordata : OUT STD_LOGIC;
                    signal txd : OUT STD_LOGIC
                 );
end component uart_1;

component niosII_system_reset_clk_0_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component niosII_system_reset_clk_0_domain_synch_module;

component niosII_system_reset_altpll_inst_c1_out_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component niosII_system_reset_altpll_inst_c1_out_domain_synch_module;

                signal altpll_inst_c1_out_reset_n :  STD_LOGIC;
                signal altpll_inst_pll_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal altpll_inst_pll_slave_read :  STD_LOGIC;
                signal altpll_inst_pll_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal altpll_inst_pll_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal altpll_inst_pll_slave_reset :  STD_LOGIC;
                signal altpll_inst_pll_slave_write :  STD_LOGIC;
                signal altpll_inst_pll_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clk_0_reset_n :  STD_LOGIC;
                signal cpu_data_master_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_data_master_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_data_master_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_data_master_byteenable_niosII_system_burst_11_upstream :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_byteenable_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal cpu_data_master_byteenable_niosII_system_burst_20_upstream :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_dbs_write_16 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal cpu_data_master_dbs_write_8 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal cpu_data_master_debugaccess :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal cpu_data_master_granted_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal cpu_data_master_irq :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_data_master_latency_counter :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal cpu_data_master_qualified_request_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal cpu_data_master_read :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register :  STD_LOGIC;
                signal cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_data_master_readdatavalid :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_11_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_13_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_14_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_15_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_16_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_17_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_18_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_1_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_20_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_21_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_3_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_4_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_5_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_6_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_7_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_8_upstream :  STD_LOGIC;
                signal cpu_data_master_requests_niosII_system_burst_9_upstream :  STD_LOGIC;
                signal cpu_data_master_waitrequest :  STD_LOGIC;
                signal cpu_data_master_write :  STD_LOGIC;
                signal cpu_data_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_instruction_master_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_instruction_master_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_granted_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal cpu_instruction_master_granted_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal cpu_instruction_master_granted_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal cpu_instruction_master_granted_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal cpu_instruction_master_granted_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal cpu_instruction_master_latency_counter :  STD_LOGIC;
                signal cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal cpu_instruction_master_read :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register :  STD_LOGIC;
                signal cpu_instruction_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal cpu_instruction_master_requests_niosII_system_burst_0_upstream :  STD_LOGIC;
                signal cpu_instruction_master_requests_niosII_system_burst_10_upstream :  STD_LOGIC;
                signal cpu_instruction_master_requests_niosII_system_burst_12_upstream :  STD_LOGIC;
                signal cpu_instruction_master_requests_niosII_system_burst_19_upstream :  STD_LOGIC;
                signal cpu_instruction_master_requests_niosII_system_burst_2_upstream :  STD_LOGIC;
                signal cpu_instruction_master_waitrequest :  STD_LOGIC;
                signal cpu_jtag_debug_module_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal cpu_jtag_debug_module_begintransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_jtag_debug_module_chipselect :  STD_LOGIC;
                signal cpu_jtag_debug_module_debugaccess :  STD_LOGIC;
                signal cpu_jtag_debug_module_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_jtag_debug_module_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_jtag_debug_module_reset_n :  STD_LOGIC;
                signal cpu_jtag_debug_module_resetrequest :  STD_LOGIC;
                signal cpu_jtag_debug_module_resetrequest_from_sa :  STD_LOGIC;
                signal cpu_jtag_debug_module_write :  STD_LOGIC;
                signal cpu_jtag_debug_module_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal d1_altpll_inst_pll_slave_end_xfer :  STD_LOGIC;
                signal d1_cpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal d1_dm9000a_inst_avalon_slave_0_end_xfer :  STD_LOGIC;
                signal d1_high_res_timer_s1_end_xfer :  STD_LOGIC;
                signal d1_jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal d1_lcd_display_control_slave_end_xfer :  STD_LOGIC;
                signal d1_led_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_memory_s1_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_0_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_10_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_11_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_12_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_13_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_14_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_15_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_16_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_17_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_18_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_19_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_1_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_20_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_21_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_2_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_3_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_4_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_5_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_6_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_7_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_8_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_burst_9_upstream_end_xfer :  STD_LOGIC;
                signal d1_niosII_system_clock_0_in_end_xfer :  STD_LOGIC;
                signal d1_sdram_s1_end_xfer :  STD_LOGIC;
                signal d1_seven_seg_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_switch_s1_end_xfer :  STD_LOGIC;
                signal d1_sys_clk_timer_s1_end_xfer :  STD_LOGIC;
                signal d1_sysid_control_slave_end_xfer :  STD_LOGIC;
                signal d1_tri_state_bridge_avalon_slave_end_xfer :  STD_LOGIC;
                signal d1_tsb_avalon_slave_end_xfer :  STD_LOGIC;
                signal d1_uart_0_s1_end_xfer :  STD_LOGIC;
                signal d1_uart_1_s1_end_xfer :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_address :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_chipselect_n :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_irq :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_irq_from_sa :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_read_n :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dm9000a_inst_avalon_slave_0_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dm9000a_inst_avalon_slave_0_reset_n :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_write_n :  STD_LOGIC;
                signal dm9000a_inst_avalon_slave_0_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal ext_flash_s1_wait_counter_eq_0 :  STD_LOGIC;
                signal high_res_timer_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal high_res_timer_s1_chipselect :  STD_LOGIC;
                signal high_res_timer_s1_irq :  STD_LOGIC;
                signal high_res_timer_s1_irq_from_sa :  STD_LOGIC;
                signal high_res_timer_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal high_res_timer_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal high_res_timer_s1_reset_n :  STD_LOGIC;
                signal high_res_timer_s1_write_n :  STD_LOGIC;
                signal high_res_timer_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal incoming_sram_IF_0_tsb_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_ENET_CMD_from_the_dm9000a_inst :  STD_LOGIC;
                signal internal_ENET_CS_N_from_the_dm9000a_inst :  STD_LOGIC;
                signal internal_ENET_RD_N_from_the_dm9000a_inst :  STD_LOGIC;
                signal internal_ENET_RST_N_from_the_dm9000a_inst :  STD_LOGIC;
                signal internal_ENET_WR_N_from_the_dm9000a_inst :  STD_LOGIC;
                signal internal_LCD_E_from_the_lcd_display :  STD_LOGIC;
                signal internal_LCD_RS_from_the_lcd_display :  STD_LOGIC;
                signal internal_LCD_RW_from_the_lcd_display :  STD_LOGIC;
                signal internal_address_to_the_ext_flash :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal internal_altpll_inst_c1_out :  STD_LOGIC;
                signal internal_coe_sram_address_from_the_sram_IF_0 :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal internal_coe_sram_chipenable_n_from_the_sram_IF_0 :  STD_LOGIC;
                signal internal_coe_sram_lowerbyte_n_from_the_sram_IF_0 :  STD_LOGIC;
                signal internal_coe_sram_outputenable_n_from_the_sram_IF_0 :  STD_LOGIC;
                signal internal_coe_sram_upperbyte_n_from_the_sram_IF_0 :  STD_LOGIC;
                signal internal_coe_sram_writeenable_n_from_the_sram_IF_0 :  STD_LOGIC;
                signal internal_locked_from_the_altpll_inst :  STD_LOGIC;
                signal internal_out_port_from_the_led_pio :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_out_port_from_the_seven_seg_pio :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_phasedone_from_the_altpll_inst :  STD_LOGIC;
                signal internal_read_n_to_the_ext_flash :  STD_LOGIC;
                signal internal_select_n_to_the_ext_flash :  STD_LOGIC;
                signal internal_txd_from_the_uart_0 :  STD_LOGIC;
                signal internal_txd_from_the_uart_1 :  STD_LOGIC;
                signal internal_write_n_to_the_ext_flash :  STD_LOGIC;
                signal internal_zs_addr_from_the_sdram :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal internal_zs_ba_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_cas_n_from_the_sdram :  STD_LOGIC;
                signal internal_zs_cke_from_the_sdram :  STD_LOGIC;
                signal internal_zs_cs_n_from_the_sdram :  STD_LOGIC;
                signal internal_zs_dqm_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_ras_n_from_the_sdram :  STD_LOGIC;
                signal internal_zs_we_n_from_the_sdram :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_address :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_chipselect :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_read_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readyfordata :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reset_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_write_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_display_control_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal lcd_display_control_slave_begintransfer :  STD_LOGIC;
                signal lcd_display_control_slave_read :  STD_LOGIC;
                signal lcd_display_control_slave_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal lcd_display_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal lcd_display_control_slave_wait_counter_eq_0 :  STD_LOGIC;
                signal lcd_display_control_slave_write :  STD_LOGIC;
                signal lcd_display_control_slave_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal led_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal led_pio_s1_chipselect :  STD_LOGIC;
                signal led_pio_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal led_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal led_pio_s1_reset_n :  STD_LOGIC;
                signal led_pio_s1_write_n :  STD_LOGIC;
                signal led_pio_s1_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal memory_s1_address :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal memory_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal memory_s1_chipselect :  STD_LOGIC;
                signal memory_s1_clken :  STD_LOGIC;
                signal memory_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal memory_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal memory_s1_reset :  STD_LOGIC;
                signal memory_s1_write :  STD_LOGIC;
                signal memory_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal module_input138 :  STD_LOGIC;
                signal module_input139 :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_0_downstream_address_to_slave :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_0_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_0_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_0_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_0_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_0_upstream_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_0_upstream_byteaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal niosII_system_burst_0_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_0_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_0_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_0_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_0_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_10_downstream_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_10_downstream_address_to_slave :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_10_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_10_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_10_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_10_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_10_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_10_upstream_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_10_upstream_byteaddress :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal niosII_system_burst_10_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_10_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_10_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_10_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_10_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_11_downstream_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_11_downstream_address_to_slave :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_11_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_11_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_11_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_11_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_11_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_11_upstream_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_11_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_11_upstream_byteaddress :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal niosII_system_burst_11_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_11_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_11_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_11_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_11_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_12_downstream_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_12_downstream_address_to_slave :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_12_downstream_arbitrationshare :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_12_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_byteenable :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_granted_ext_flash_s1 :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_12_downstream_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1 :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_12_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_requests_ext_flash_s1 :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_12_upstream_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_12_upstream_byteaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_12_upstream_byteenable :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_12_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_12_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_12_upstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_13_downstream_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_13_downstream_address_to_slave :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_13_downstream_arbitrationshare :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_13_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_byteenable :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_granted_ext_flash_s1 :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_13_downstream_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1 :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_13_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_requests_ext_flash_s1 :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_13_upstream_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_13_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_13_upstream_byteaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_13_upstream_byteenable :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_13_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_13_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_13_upstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_14_downstream_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_14_downstream_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_14_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_14_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_14_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1 :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_14_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_14_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_14_upstream_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_14_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_14_upstream_byteaddress :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_14_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_14_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_14_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_14_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_14_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_15_downstream_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_downstream_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_15_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_15_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_granted_high_res_timer_s1 :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_nativeaddress :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1 :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_15_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_requests_high_res_timer_s1 :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_15_upstream_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_15_upstream_byteaddress :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_15_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_15_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_15_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_15_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_15_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_16_downstream_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_16_downstream_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_16_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_16_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_16_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0 :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_16_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_16_upstream_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_16_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_16_upstream_byteaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_16_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_16_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_16_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_16_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_16_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_17_downstream_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_downstream_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_17_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_17_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_granted_uart_0_s1 :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_nativeaddress :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_downstream_qualified_request_uart_0_s1 :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_read_data_valid_uart_0_s1 :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_17_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_requests_uart_0_s1 :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_17_upstream_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_17_upstream_byteaddress :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_17_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_17_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_17_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_17_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_17_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_18_downstream_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_downstream_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_18_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_18_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_granted_uart_1_s1 :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_nativeaddress :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_downstream_qualified_request_uart_1_s1 :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_read_data_valid_uart_1_s1 :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_18_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_requests_uart_1_s1 :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_18_upstream_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_18_upstream_byteaddress :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_18_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_18_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_18_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_18_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_18_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_19_downstream_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_19_downstream_address_to_slave :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_19_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_19_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_19_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_granted_sram_IF_0_tsb :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_19_downstream_nativeaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_19_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_requests_sram_IF_0_tsb :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_19_upstream_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_19_upstream_byteaddress :  STD_LOGIC_VECTOR (19 DOWNTO 0);
                signal niosII_system_burst_19_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_19_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_19_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_19_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_19_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_1_downstream_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_1_downstream_address_to_slave :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_1_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_1_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_1_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_1_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_1_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_1_upstream_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_1_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_1_upstream_byteaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal niosII_system_burst_1_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_1_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_1_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_1_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_1_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_20_downstream_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_20_downstream_address_to_slave :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_20_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_20_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_20_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_granted_sram_IF_0_tsb :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_20_downstream_nativeaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_20_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_requests_sram_IF_0_tsb :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_20_upstream_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_20_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_20_upstream_byteaddress :  STD_LOGIC_VECTOR (19 DOWNTO 0);
                signal niosII_system_burst_20_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_20_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_20_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_20_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_20_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_21_downstream_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_downstream_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_nativeaddress :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_21_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_21_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_21_upstream_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_upstream_byteaddress :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_21_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_21_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_21_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_21_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_21_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_2_downstream_address :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_2_downstream_address_to_slave :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_2_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_2_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_2_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_granted_memory_s1 :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_nativeaddress :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_2_downstream_qualified_request_memory_s1 :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_read_data_valid_memory_s1 :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_2_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_requests_memory_s1 :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_2_upstream_address :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_2_upstream_byteaddress :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_2_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_2_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_2_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_2_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_2_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_3_downstream_address :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_3_downstream_address_to_slave :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_3_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_3_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_3_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_granted_memory_s1 :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_nativeaddress :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_3_downstream_qualified_request_memory_s1 :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_read_data_valid_memory_s1 :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_3_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_requests_memory_s1 :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_3_upstream_address :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_3_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_3_upstream_byteaddress :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_3_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_3_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_3_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_3_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_3_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_4_downstream_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_4_downstream_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_4_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_4_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_4_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_granted_sysid_control_slave :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_4_downstream_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_4_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_requests_sysid_control_slave :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_4_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_4_upstream_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_4_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_4_upstream_byteaddress :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_4_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_4_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_4_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_4_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_4_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_5_downstream_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_downstream_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_5_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_5_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_nativeaddress :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1 :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_5_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_5_upstream_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_5_upstream_byteaddress :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_5_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_5_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_5_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_5_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_5_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_6_downstream_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_6_downstream_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_6_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_6_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_6_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_6_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_6_upstream_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_system_burst_6_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_6_upstream_byteaddress :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal niosII_system_burst_6_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_6_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_6_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_6_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_6_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_7_downstream_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_7_downstream_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_7_downstream_arbitrationshare :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_7_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_byteenable :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_granted_lcd_display_control_slave :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_7_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_requests_lcd_display_control_slave :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_7_upstream_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_7_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_7_upstream_byteaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_7_upstream_byteenable :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_7_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_7_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_7_upstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_8_downstream_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_8_downstream_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_8_downstream_arbitrationshare :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_8_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_byteenable :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_granted_led_pio_s1 :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_8_downstream_qualified_request_led_pio_s1 :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_read_data_valid_led_pio_s1 :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_8_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_requests_led_pio_s1 :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_8_upstream_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_8_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_8_upstream_byteaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_8_upstream_byteenable :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_8_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_8_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_8_upstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_9_downstream_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_9_downstream_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_9_downstream_arbitrationshare :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_system_burst_9_downstream_burstcount :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_byteenable :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_granted_switch_s1 :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_latency_counter :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_9_downstream_qualified_request_switch_s1 :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_read :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_read_data_valid_switch_s1 :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_9_downstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_requests_switch_s1 :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_reset_n :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_write :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_9_upstream_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_9_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_burst_9_upstream_byteaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_burst_9_upstream_byteenable :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_read :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_9_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_9_upstream_readdatavalid :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_waitrequest :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_write :  STD_LOGIC;
                signal niosII_system_burst_9_upstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_clock_0_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_clock_0_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_clock_0_in_endofpacket :  STD_LOGIC;
                signal niosII_system_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_system_clock_0_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_clock_0_in_read :  STD_LOGIC;
                signal niosII_system_clock_0_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_clock_0_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_clock_0_in_reset_n :  STD_LOGIC;
                signal niosII_system_clock_0_in_waitrequest :  STD_LOGIC;
                signal niosII_system_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_system_clock_0_in_write :  STD_LOGIC;
                signal niosII_system_clock_0_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_clock_0_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_clock_0_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_system_clock_0_out_endofpacket :  STD_LOGIC;
                signal niosII_system_clock_0_out_granted_altpll_inst_pll_slave :  STD_LOGIC;
                signal niosII_system_clock_0_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave :  STD_LOGIC;
                signal niosII_system_clock_0_out_read :  STD_LOGIC;
                signal niosII_system_clock_0_out_read_data_valid_altpll_inst_pll_slave :  STD_LOGIC;
                signal niosII_system_clock_0_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_clock_0_out_requests_altpll_inst_pll_slave :  STD_LOGIC;
                signal niosII_system_clock_0_out_reset_n :  STD_LOGIC;
                signal niosII_system_clock_0_out_waitrequest :  STD_LOGIC;
                signal niosII_system_clock_0_out_write :  STD_LOGIC;
                signal niosII_system_clock_0_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal out_clk_altpll_inst_c0 :  STD_LOGIC;
                signal out_clk_altpll_inst_c1 :  STD_LOGIC;
                signal out_clk_altpll_inst_c2 :  STD_LOGIC;
                signal reset_n_sources :  STD_LOGIC;
                signal sdram_s1_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal sdram_s1_byteenable_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_s1_chipselect :  STD_LOGIC;
                signal sdram_s1_read_n :  STD_LOGIC;
                signal sdram_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sdram_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sdram_s1_readdatavalid :  STD_LOGIC;
                signal sdram_s1_reset_n :  STD_LOGIC;
                signal sdram_s1_waitrequest :  STD_LOGIC;
                signal sdram_s1_waitrequest_from_sa :  STD_LOGIC;
                signal sdram_s1_write_n :  STD_LOGIC;
                signal sdram_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal seven_seg_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal seven_seg_pio_s1_chipselect :  STD_LOGIC;
                signal seven_seg_pio_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal seven_seg_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal seven_seg_pio_s1_reset_n :  STD_LOGIC;
                signal seven_seg_pio_s1_write_n :  STD_LOGIC;
                signal seven_seg_pio_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sram_IF_0_tsb_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal sram_IF_0_tsb_byteenable_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sram_IF_0_tsb_chipselect_n :  STD_LOGIC;
                signal sram_IF_0_tsb_outputenable_n :  STD_LOGIC;
                signal sram_IF_0_tsb_write_n :  STD_LOGIC;
                signal switch_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal switch_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal switch_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal switch_s1_reset_n :  STD_LOGIC;
                signal sys_clk_timer_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sys_clk_timer_s1_chipselect :  STD_LOGIC;
                signal sys_clk_timer_s1_irq :  STD_LOGIC;
                signal sys_clk_timer_s1_irq_from_sa :  STD_LOGIC;
                signal sys_clk_timer_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sys_clk_timer_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sys_clk_timer_s1_reset_n :  STD_LOGIC;
                signal sys_clk_timer_s1_write_n :  STD_LOGIC;
                signal sys_clk_timer_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sysid_control_slave_address :  STD_LOGIC;
                signal sysid_control_slave_clock :  STD_LOGIC;
                signal sysid_control_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_reset_n :  STD_LOGIC;
                signal uart_0_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal uart_0_s1_begintransfer :  STD_LOGIC;
                signal uart_0_s1_chipselect :  STD_LOGIC;
                signal uart_0_s1_dataavailable :  STD_LOGIC;
                signal uart_0_s1_dataavailable_from_sa :  STD_LOGIC;
                signal uart_0_s1_irq :  STD_LOGIC;
                signal uart_0_s1_irq_from_sa :  STD_LOGIC;
                signal uart_0_s1_read_n :  STD_LOGIC;
                signal uart_0_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal uart_0_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal uart_0_s1_readyfordata :  STD_LOGIC;
                signal uart_0_s1_readyfordata_from_sa :  STD_LOGIC;
                signal uart_0_s1_reset_n :  STD_LOGIC;
                signal uart_0_s1_write_n :  STD_LOGIC;
                signal uart_0_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal uart_1_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal uart_1_s1_begintransfer :  STD_LOGIC;
                signal uart_1_s1_chipselect :  STD_LOGIC;
                signal uart_1_s1_dataavailable :  STD_LOGIC;
                signal uart_1_s1_dataavailable_from_sa :  STD_LOGIC;
                signal uart_1_s1_irq :  STD_LOGIC;
                signal uart_1_s1_irq_from_sa :  STD_LOGIC;
                signal uart_1_s1_read_n :  STD_LOGIC;
                signal uart_1_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal uart_1_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal uart_1_s1_readyfordata :  STD_LOGIC;
                signal uart_1_s1_readyfordata_from_sa :  STD_LOGIC;
                signal uart_1_s1_reset_n :  STD_LOGIC;
                signal uart_1_s1_write_n :  STD_LOGIC;
                signal uart_1_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);

begin

  --the_altpll_inst_pll_slave, which is an e_instance
  the_altpll_inst_pll_slave : altpll_inst_pll_slave_arbitrator
    port map(
      altpll_inst_pll_slave_address => altpll_inst_pll_slave_address,
      altpll_inst_pll_slave_read => altpll_inst_pll_slave_read,
      altpll_inst_pll_slave_readdata_from_sa => altpll_inst_pll_slave_readdata_from_sa,
      altpll_inst_pll_slave_reset => altpll_inst_pll_slave_reset,
      altpll_inst_pll_slave_write => altpll_inst_pll_slave_write,
      altpll_inst_pll_slave_writedata => altpll_inst_pll_slave_writedata,
      d1_altpll_inst_pll_slave_end_xfer => d1_altpll_inst_pll_slave_end_xfer,
      niosII_system_clock_0_out_granted_altpll_inst_pll_slave => niosII_system_clock_0_out_granted_altpll_inst_pll_slave,
      niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave => niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave,
      niosII_system_clock_0_out_read_data_valid_altpll_inst_pll_slave => niosII_system_clock_0_out_read_data_valid_altpll_inst_pll_slave,
      niosII_system_clock_0_out_requests_altpll_inst_pll_slave => niosII_system_clock_0_out_requests_altpll_inst_pll_slave,
      altpll_inst_pll_slave_readdata => altpll_inst_pll_slave_readdata,
      clk => clk_0,
      niosII_system_clock_0_out_address_to_slave => niosII_system_clock_0_out_address_to_slave,
      niosII_system_clock_0_out_read => niosII_system_clock_0_out_read,
      niosII_system_clock_0_out_write => niosII_system_clock_0_out_write,
      niosII_system_clock_0_out_writedata => niosII_system_clock_0_out_writedata,
      reset_n => clk_0_reset_n
    );


  --altpll_inst_c0_out out_clk assignment, which is an e_assign
  altpll_inst_c0_out <= out_clk_altpll_inst_c0;
  --altpll_inst_c1_out out_clk assignment, which is an e_assign
  internal_altpll_inst_c1_out <= out_clk_altpll_inst_c1;
  --altpll_inst_c2_out out_clk assignment, which is an e_assign
  altpll_inst_c2_out <= out_clk_altpll_inst_c2;
  --the_altpll_inst, which is an e_ptf_instance
  the_altpll_inst : altpll_inst
    port map(
      c0 => out_clk_altpll_inst_c0,
      c1 => out_clk_altpll_inst_c1,
      c2 => out_clk_altpll_inst_c2,
      locked => internal_locked_from_the_altpll_inst,
      phasedone => internal_phasedone_from_the_altpll_inst,
      readdata => altpll_inst_pll_slave_readdata,
      address => altpll_inst_pll_slave_address,
      clk => clk_0,
      read => altpll_inst_pll_slave_read,
      reset => altpll_inst_pll_slave_reset,
      write => altpll_inst_pll_slave_write,
      writedata => altpll_inst_pll_slave_writedata
    );


  --the_cpu_jtag_debug_module, which is an e_instance
  the_cpu_jtag_debug_module : cpu_jtag_debug_module_arbitrator
    port map(
      cpu_jtag_debug_module_address => cpu_jtag_debug_module_address,
      cpu_jtag_debug_module_begintransfer => cpu_jtag_debug_module_begintransfer,
      cpu_jtag_debug_module_byteenable => cpu_jtag_debug_module_byteenable,
      cpu_jtag_debug_module_chipselect => cpu_jtag_debug_module_chipselect,
      cpu_jtag_debug_module_debugaccess => cpu_jtag_debug_module_debugaccess,
      cpu_jtag_debug_module_readdata_from_sa => cpu_jtag_debug_module_readdata_from_sa,
      cpu_jtag_debug_module_reset_n => cpu_jtag_debug_module_reset_n,
      cpu_jtag_debug_module_resetrequest_from_sa => cpu_jtag_debug_module_resetrequest_from_sa,
      cpu_jtag_debug_module_write => cpu_jtag_debug_module_write,
      cpu_jtag_debug_module_writedata => cpu_jtag_debug_module_writedata,
      d1_cpu_jtag_debug_module_end_xfer => d1_cpu_jtag_debug_module_end_xfer,
      niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module => niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module,
      niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module => niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module,
      niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module => niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module,
      niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module => niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module,
      niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module => niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module,
      niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module => niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module,
      niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module => niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module,
      niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module => niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module,
      clk => internal_altpll_inst_c1_out,
      cpu_jtag_debug_module_readdata => cpu_jtag_debug_module_readdata,
      cpu_jtag_debug_module_resetrequest => cpu_jtag_debug_module_resetrequest,
      niosII_system_burst_0_downstream_address_to_slave => niosII_system_burst_0_downstream_address_to_slave,
      niosII_system_burst_0_downstream_arbitrationshare => niosII_system_burst_0_downstream_arbitrationshare,
      niosII_system_burst_0_downstream_burstcount => niosII_system_burst_0_downstream_burstcount,
      niosII_system_burst_0_downstream_byteenable => niosII_system_burst_0_downstream_byteenable,
      niosII_system_burst_0_downstream_debugaccess => niosII_system_burst_0_downstream_debugaccess,
      niosII_system_burst_0_downstream_latency_counter => niosII_system_burst_0_downstream_latency_counter,
      niosII_system_burst_0_downstream_read => niosII_system_burst_0_downstream_read,
      niosII_system_burst_0_downstream_write => niosII_system_burst_0_downstream_write,
      niosII_system_burst_0_downstream_writedata => niosII_system_burst_0_downstream_writedata,
      niosII_system_burst_1_downstream_address_to_slave => niosII_system_burst_1_downstream_address_to_slave,
      niosII_system_burst_1_downstream_arbitrationshare => niosII_system_burst_1_downstream_arbitrationshare,
      niosII_system_burst_1_downstream_burstcount => niosII_system_burst_1_downstream_burstcount,
      niosII_system_burst_1_downstream_byteenable => niosII_system_burst_1_downstream_byteenable,
      niosII_system_burst_1_downstream_debugaccess => niosII_system_burst_1_downstream_debugaccess,
      niosII_system_burst_1_downstream_latency_counter => niosII_system_burst_1_downstream_latency_counter,
      niosII_system_burst_1_downstream_read => niosII_system_burst_1_downstream_read,
      niosII_system_burst_1_downstream_write => niosII_system_burst_1_downstream_write,
      niosII_system_burst_1_downstream_writedata => niosII_system_burst_1_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_cpu_data_master, which is an e_instance
  the_cpu_data_master : cpu_data_master_arbitrator
    port map(
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_dbs_address => cpu_data_master_dbs_address,
      cpu_data_master_dbs_write_16 => cpu_data_master_dbs_write_16,
      cpu_data_master_dbs_write_8 => cpu_data_master_dbs_write_8,
      cpu_data_master_irq => cpu_data_master_irq,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_readdata => cpu_data_master_readdata,
      cpu_data_master_readdatavalid => cpu_data_master_readdatavalid,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address => cpu_data_master_address,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_byteenable_niosII_system_burst_11_upstream => cpu_data_master_byteenable_niosII_system_burst_11_upstream,
      cpu_data_master_byteenable_niosII_system_burst_13_upstream => cpu_data_master_byteenable_niosII_system_burst_13_upstream,
      cpu_data_master_byteenable_niosII_system_burst_20_upstream => cpu_data_master_byteenable_niosII_system_burst_20_upstream,
      cpu_data_master_granted_niosII_system_burst_11_upstream => cpu_data_master_granted_niosII_system_burst_11_upstream,
      cpu_data_master_granted_niosII_system_burst_13_upstream => cpu_data_master_granted_niosII_system_burst_13_upstream,
      cpu_data_master_granted_niosII_system_burst_14_upstream => cpu_data_master_granted_niosII_system_burst_14_upstream,
      cpu_data_master_granted_niosII_system_burst_15_upstream => cpu_data_master_granted_niosII_system_burst_15_upstream,
      cpu_data_master_granted_niosII_system_burst_16_upstream => cpu_data_master_granted_niosII_system_burst_16_upstream,
      cpu_data_master_granted_niosII_system_burst_17_upstream => cpu_data_master_granted_niosII_system_burst_17_upstream,
      cpu_data_master_granted_niosII_system_burst_18_upstream => cpu_data_master_granted_niosII_system_burst_18_upstream,
      cpu_data_master_granted_niosII_system_burst_1_upstream => cpu_data_master_granted_niosII_system_burst_1_upstream,
      cpu_data_master_granted_niosII_system_burst_20_upstream => cpu_data_master_granted_niosII_system_burst_20_upstream,
      cpu_data_master_granted_niosII_system_burst_21_upstream => cpu_data_master_granted_niosII_system_burst_21_upstream,
      cpu_data_master_granted_niosII_system_burst_3_upstream => cpu_data_master_granted_niosII_system_burst_3_upstream,
      cpu_data_master_granted_niosII_system_burst_4_upstream => cpu_data_master_granted_niosII_system_burst_4_upstream,
      cpu_data_master_granted_niosII_system_burst_5_upstream => cpu_data_master_granted_niosII_system_burst_5_upstream,
      cpu_data_master_granted_niosII_system_burst_6_upstream => cpu_data_master_granted_niosII_system_burst_6_upstream,
      cpu_data_master_granted_niosII_system_burst_7_upstream => cpu_data_master_granted_niosII_system_burst_7_upstream,
      cpu_data_master_granted_niosII_system_burst_8_upstream => cpu_data_master_granted_niosII_system_burst_8_upstream,
      cpu_data_master_granted_niosII_system_burst_9_upstream => cpu_data_master_granted_niosII_system_burst_9_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_11_upstream => cpu_data_master_qualified_request_niosII_system_burst_11_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_13_upstream => cpu_data_master_qualified_request_niosII_system_burst_13_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_14_upstream => cpu_data_master_qualified_request_niosII_system_burst_14_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_15_upstream => cpu_data_master_qualified_request_niosII_system_burst_15_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_16_upstream => cpu_data_master_qualified_request_niosII_system_burst_16_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_17_upstream => cpu_data_master_qualified_request_niosII_system_burst_17_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_18_upstream => cpu_data_master_qualified_request_niosII_system_burst_18_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_1_upstream => cpu_data_master_qualified_request_niosII_system_burst_1_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_20_upstream => cpu_data_master_qualified_request_niosII_system_burst_20_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_21_upstream => cpu_data_master_qualified_request_niosII_system_burst_21_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_3_upstream => cpu_data_master_qualified_request_niosII_system_burst_3_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_4_upstream => cpu_data_master_qualified_request_niosII_system_burst_4_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_5_upstream => cpu_data_master_qualified_request_niosII_system_burst_5_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_6_upstream => cpu_data_master_qualified_request_niosII_system_burst_6_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_7_upstream => cpu_data_master_qualified_request_niosII_system_burst_7_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_8_upstream => cpu_data_master_qualified_request_niosII_system_burst_8_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_9_upstream => cpu_data_master_qualified_request_niosII_system_burst_9_upstream,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_11_upstream => cpu_data_master_requests_niosII_system_burst_11_upstream,
      cpu_data_master_requests_niosII_system_burst_13_upstream => cpu_data_master_requests_niosII_system_burst_13_upstream,
      cpu_data_master_requests_niosII_system_burst_14_upstream => cpu_data_master_requests_niosII_system_burst_14_upstream,
      cpu_data_master_requests_niosII_system_burst_15_upstream => cpu_data_master_requests_niosII_system_burst_15_upstream,
      cpu_data_master_requests_niosII_system_burst_16_upstream => cpu_data_master_requests_niosII_system_burst_16_upstream,
      cpu_data_master_requests_niosII_system_burst_17_upstream => cpu_data_master_requests_niosII_system_burst_17_upstream,
      cpu_data_master_requests_niosII_system_burst_18_upstream => cpu_data_master_requests_niosII_system_burst_18_upstream,
      cpu_data_master_requests_niosII_system_burst_1_upstream => cpu_data_master_requests_niosII_system_burst_1_upstream,
      cpu_data_master_requests_niosII_system_burst_20_upstream => cpu_data_master_requests_niosII_system_burst_20_upstream,
      cpu_data_master_requests_niosII_system_burst_21_upstream => cpu_data_master_requests_niosII_system_burst_21_upstream,
      cpu_data_master_requests_niosII_system_burst_3_upstream => cpu_data_master_requests_niosII_system_burst_3_upstream,
      cpu_data_master_requests_niosII_system_burst_4_upstream => cpu_data_master_requests_niosII_system_burst_4_upstream,
      cpu_data_master_requests_niosII_system_burst_5_upstream => cpu_data_master_requests_niosII_system_burst_5_upstream,
      cpu_data_master_requests_niosII_system_burst_6_upstream => cpu_data_master_requests_niosII_system_burst_6_upstream,
      cpu_data_master_requests_niosII_system_burst_7_upstream => cpu_data_master_requests_niosII_system_burst_7_upstream,
      cpu_data_master_requests_niosII_system_burst_8_upstream => cpu_data_master_requests_niosII_system_burst_8_upstream,
      cpu_data_master_requests_niosII_system_burst_9_upstream => cpu_data_master_requests_niosII_system_burst_9_upstream,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      d1_niosII_system_burst_11_upstream_end_xfer => d1_niosII_system_burst_11_upstream_end_xfer,
      d1_niosII_system_burst_13_upstream_end_xfer => d1_niosII_system_burst_13_upstream_end_xfer,
      d1_niosII_system_burst_14_upstream_end_xfer => d1_niosII_system_burst_14_upstream_end_xfer,
      d1_niosII_system_burst_15_upstream_end_xfer => d1_niosII_system_burst_15_upstream_end_xfer,
      d1_niosII_system_burst_16_upstream_end_xfer => d1_niosII_system_burst_16_upstream_end_xfer,
      d1_niosII_system_burst_17_upstream_end_xfer => d1_niosII_system_burst_17_upstream_end_xfer,
      d1_niosII_system_burst_18_upstream_end_xfer => d1_niosII_system_burst_18_upstream_end_xfer,
      d1_niosII_system_burst_1_upstream_end_xfer => d1_niosII_system_burst_1_upstream_end_xfer,
      d1_niosII_system_burst_20_upstream_end_xfer => d1_niosII_system_burst_20_upstream_end_xfer,
      d1_niosII_system_burst_21_upstream_end_xfer => d1_niosII_system_burst_21_upstream_end_xfer,
      d1_niosII_system_burst_3_upstream_end_xfer => d1_niosII_system_burst_3_upstream_end_xfer,
      d1_niosII_system_burst_4_upstream_end_xfer => d1_niosII_system_burst_4_upstream_end_xfer,
      d1_niosII_system_burst_5_upstream_end_xfer => d1_niosII_system_burst_5_upstream_end_xfer,
      d1_niosII_system_burst_6_upstream_end_xfer => d1_niosII_system_burst_6_upstream_end_xfer,
      d1_niosII_system_burst_7_upstream_end_xfer => d1_niosII_system_burst_7_upstream_end_xfer,
      d1_niosII_system_burst_8_upstream_end_xfer => d1_niosII_system_burst_8_upstream_end_xfer,
      d1_niosII_system_burst_9_upstream_end_xfer => d1_niosII_system_burst_9_upstream_end_xfer,
      dm9000a_inst_avalon_slave_0_irq_from_sa => dm9000a_inst_avalon_slave_0_irq_from_sa,
      high_res_timer_s1_irq_from_sa => high_res_timer_s1_irq_from_sa,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      niosII_system_burst_11_upstream_readdata_from_sa => niosII_system_burst_11_upstream_readdata_from_sa,
      niosII_system_burst_11_upstream_waitrequest_from_sa => niosII_system_burst_11_upstream_waitrequest_from_sa,
      niosII_system_burst_13_upstream_readdata_from_sa => niosII_system_burst_13_upstream_readdata_from_sa,
      niosII_system_burst_13_upstream_waitrequest_from_sa => niosII_system_burst_13_upstream_waitrequest_from_sa,
      niosII_system_burst_14_upstream_readdata_from_sa => niosII_system_burst_14_upstream_readdata_from_sa,
      niosII_system_burst_14_upstream_waitrequest_from_sa => niosII_system_burst_14_upstream_waitrequest_from_sa,
      niosII_system_burst_15_upstream_readdata_from_sa => niosII_system_burst_15_upstream_readdata_from_sa,
      niosII_system_burst_15_upstream_waitrequest_from_sa => niosII_system_burst_15_upstream_waitrequest_from_sa,
      niosII_system_burst_16_upstream_readdata_from_sa => niosII_system_burst_16_upstream_readdata_from_sa,
      niosII_system_burst_16_upstream_waitrequest_from_sa => niosII_system_burst_16_upstream_waitrequest_from_sa,
      niosII_system_burst_17_upstream_readdata_from_sa => niosII_system_burst_17_upstream_readdata_from_sa,
      niosII_system_burst_17_upstream_waitrequest_from_sa => niosII_system_burst_17_upstream_waitrequest_from_sa,
      niosII_system_burst_18_upstream_readdata_from_sa => niosII_system_burst_18_upstream_readdata_from_sa,
      niosII_system_burst_18_upstream_waitrequest_from_sa => niosII_system_burst_18_upstream_waitrequest_from_sa,
      niosII_system_burst_1_upstream_readdata_from_sa => niosII_system_burst_1_upstream_readdata_from_sa,
      niosII_system_burst_1_upstream_waitrequest_from_sa => niosII_system_burst_1_upstream_waitrequest_from_sa,
      niosII_system_burst_20_upstream_readdata_from_sa => niosII_system_burst_20_upstream_readdata_from_sa,
      niosII_system_burst_20_upstream_waitrequest_from_sa => niosII_system_burst_20_upstream_waitrequest_from_sa,
      niosII_system_burst_21_upstream_readdata_from_sa => niosII_system_burst_21_upstream_readdata_from_sa,
      niosII_system_burst_21_upstream_waitrequest_from_sa => niosII_system_burst_21_upstream_waitrequest_from_sa,
      niosII_system_burst_3_upstream_readdata_from_sa => niosII_system_burst_3_upstream_readdata_from_sa,
      niosII_system_burst_3_upstream_waitrequest_from_sa => niosII_system_burst_3_upstream_waitrequest_from_sa,
      niosII_system_burst_4_upstream_readdata_from_sa => niosII_system_burst_4_upstream_readdata_from_sa,
      niosII_system_burst_4_upstream_waitrequest_from_sa => niosII_system_burst_4_upstream_waitrequest_from_sa,
      niosII_system_burst_5_upstream_readdata_from_sa => niosII_system_burst_5_upstream_readdata_from_sa,
      niosII_system_burst_5_upstream_waitrequest_from_sa => niosII_system_burst_5_upstream_waitrequest_from_sa,
      niosII_system_burst_6_upstream_readdata_from_sa => niosII_system_burst_6_upstream_readdata_from_sa,
      niosII_system_burst_6_upstream_waitrequest_from_sa => niosII_system_burst_6_upstream_waitrequest_from_sa,
      niosII_system_burst_7_upstream_readdata_from_sa => niosII_system_burst_7_upstream_readdata_from_sa,
      niosII_system_burst_7_upstream_waitrequest_from_sa => niosII_system_burst_7_upstream_waitrequest_from_sa,
      niosII_system_burst_8_upstream_readdata_from_sa => niosII_system_burst_8_upstream_readdata_from_sa,
      niosII_system_burst_8_upstream_waitrequest_from_sa => niosII_system_burst_8_upstream_waitrequest_from_sa,
      niosII_system_burst_9_upstream_readdata_from_sa => niosII_system_burst_9_upstream_readdata_from_sa,
      niosII_system_burst_9_upstream_waitrequest_from_sa => niosII_system_burst_9_upstream_waitrequest_from_sa,
      reset_n => altpll_inst_c1_out_reset_n,
      sys_clk_timer_s1_irq_from_sa => sys_clk_timer_s1_irq_from_sa,
      uart_0_s1_irq_from_sa => uart_0_s1_irq_from_sa,
      uart_1_s1_irq_from_sa => uart_1_s1_irq_from_sa
    );


  --the_cpu_instruction_master, which is an e_instance
  the_cpu_instruction_master : cpu_instruction_master_arbitrator
    port map(
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_dbs_address => cpu_instruction_master_dbs_address,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_readdata => cpu_instruction_master_readdata,
      cpu_instruction_master_readdatavalid => cpu_instruction_master_readdatavalid,
      cpu_instruction_master_waitrequest => cpu_instruction_master_waitrequest,
      clk => internal_altpll_inst_c1_out,
      cpu_instruction_master_address => cpu_instruction_master_address,
      cpu_instruction_master_burstcount => cpu_instruction_master_burstcount,
      cpu_instruction_master_granted_niosII_system_burst_0_upstream => cpu_instruction_master_granted_niosII_system_burst_0_upstream,
      cpu_instruction_master_granted_niosII_system_burst_10_upstream => cpu_instruction_master_granted_niosII_system_burst_10_upstream,
      cpu_instruction_master_granted_niosII_system_burst_12_upstream => cpu_instruction_master_granted_niosII_system_burst_12_upstream,
      cpu_instruction_master_granted_niosII_system_burst_19_upstream => cpu_instruction_master_granted_niosII_system_burst_19_upstream,
      cpu_instruction_master_granted_niosII_system_burst_2_upstream => cpu_instruction_master_granted_niosII_system_burst_2_upstream,
      cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream => cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream,
      cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream => cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream,
      cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream => cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream,
      cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream => cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream,
      cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream => cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream => cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream => cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream => cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream => cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream => cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register,
      cpu_instruction_master_requests_niosII_system_burst_0_upstream => cpu_instruction_master_requests_niosII_system_burst_0_upstream,
      cpu_instruction_master_requests_niosII_system_burst_10_upstream => cpu_instruction_master_requests_niosII_system_burst_10_upstream,
      cpu_instruction_master_requests_niosII_system_burst_12_upstream => cpu_instruction_master_requests_niosII_system_burst_12_upstream,
      cpu_instruction_master_requests_niosII_system_burst_19_upstream => cpu_instruction_master_requests_niosII_system_burst_19_upstream,
      cpu_instruction_master_requests_niosII_system_burst_2_upstream => cpu_instruction_master_requests_niosII_system_burst_2_upstream,
      d1_niosII_system_burst_0_upstream_end_xfer => d1_niosII_system_burst_0_upstream_end_xfer,
      d1_niosII_system_burst_10_upstream_end_xfer => d1_niosII_system_burst_10_upstream_end_xfer,
      d1_niosII_system_burst_12_upstream_end_xfer => d1_niosII_system_burst_12_upstream_end_xfer,
      d1_niosII_system_burst_19_upstream_end_xfer => d1_niosII_system_burst_19_upstream_end_xfer,
      d1_niosII_system_burst_2_upstream_end_xfer => d1_niosII_system_burst_2_upstream_end_xfer,
      niosII_system_burst_0_upstream_readdata_from_sa => niosII_system_burst_0_upstream_readdata_from_sa,
      niosII_system_burst_0_upstream_waitrequest_from_sa => niosII_system_burst_0_upstream_waitrequest_from_sa,
      niosII_system_burst_10_upstream_readdata_from_sa => niosII_system_burst_10_upstream_readdata_from_sa,
      niosII_system_burst_10_upstream_waitrequest_from_sa => niosII_system_burst_10_upstream_waitrequest_from_sa,
      niosII_system_burst_12_upstream_readdata_from_sa => niosII_system_burst_12_upstream_readdata_from_sa,
      niosII_system_burst_12_upstream_waitrequest_from_sa => niosII_system_burst_12_upstream_waitrequest_from_sa,
      niosII_system_burst_19_upstream_readdata_from_sa => niosII_system_burst_19_upstream_readdata_from_sa,
      niosII_system_burst_19_upstream_waitrequest_from_sa => niosII_system_burst_19_upstream_waitrequest_from_sa,
      niosII_system_burst_2_upstream_readdata_from_sa => niosII_system_burst_2_upstream_readdata_from_sa,
      niosII_system_burst_2_upstream_waitrequest_from_sa => niosII_system_burst_2_upstream_waitrequest_from_sa,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_cpu, which is an e_ptf_instance
  the_cpu : cpu
    port map(
      d_address => cpu_data_master_address,
      d_burstcount => cpu_data_master_burstcount,
      d_byteenable => cpu_data_master_byteenable,
      d_read => cpu_data_master_read,
      d_write => cpu_data_master_write,
      d_writedata => cpu_data_master_writedata,
      i_address => cpu_instruction_master_address,
      i_burstcount => cpu_instruction_master_burstcount,
      i_read => cpu_instruction_master_read,
      jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,
      jtag_debug_module_readdata => cpu_jtag_debug_module_readdata,
      jtag_debug_module_resetrequest => cpu_jtag_debug_module_resetrequest,
      clk => internal_altpll_inst_c1_out,
      d_irq => cpu_data_master_irq,
      d_readdata => cpu_data_master_readdata,
      d_readdatavalid => cpu_data_master_readdatavalid,
      d_waitrequest => cpu_data_master_waitrequest,
      i_readdata => cpu_instruction_master_readdata,
      i_readdatavalid => cpu_instruction_master_readdatavalid,
      i_waitrequest => cpu_instruction_master_waitrequest,
      jtag_debug_module_address => cpu_jtag_debug_module_address,
      jtag_debug_module_begintransfer => cpu_jtag_debug_module_begintransfer,
      jtag_debug_module_byteenable => cpu_jtag_debug_module_byteenable,
      jtag_debug_module_debugaccess => cpu_jtag_debug_module_debugaccess,
      jtag_debug_module_select => cpu_jtag_debug_module_chipselect,
      jtag_debug_module_write => cpu_jtag_debug_module_write,
      jtag_debug_module_writedata => cpu_jtag_debug_module_writedata,
      reset_n => cpu_jtag_debug_module_reset_n
    );


  --the_dm9000a_inst_avalon_slave_0, which is an e_instance
  the_dm9000a_inst_avalon_slave_0 : dm9000a_inst_avalon_slave_0_arbitrator
    port map(
      d1_dm9000a_inst_avalon_slave_0_end_xfer => d1_dm9000a_inst_avalon_slave_0_end_xfer,
      dm9000a_inst_avalon_slave_0_address => dm9000a_inst_avalon_slave_0_address,
      dm9000a_inst_avalon_slave_0_chipselect_n => dm9000a_inst_avalon_slave_0_chipselect_n,
      dm9000a_inst_avalon_slave_0_irq_from_sa => dm9000a_inst_avalon_slave_0_irq_from_sa,
      dm9000a_inst_avalon_slave_0_read_n => dm9000a_inst_avalon_slave_0_read_n,
      dm9000a_inst_avalon_slave_0_readdata_from_sa => dm9000a_inst_avalon_slave_0_readdata_from_sa,
      dm9000a_inst_avalon_slave_0_reset_n => dm9000a_inst_avalon_slave_0_reset_n,
      dm9000a_inst_avalon_slave_0_write_n => dm9000a_inst_avalon_slave_0_write_n,
      dm9000a_inst_avalon_slave_0_writedata => dm9000a_inst_avalon_slave_0_writedata,
      niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 => niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0,
      niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 => niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0,
      niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0 => niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0,
      niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 => niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0,
      clk => internal_altpll_inst_c1_out,
      dm9000a_inst_avalon_slave_0_irq => dm9000a_inst_avalon_slave_0_irq,
      dm9000a_inst_avalon_slave_0_readdata => dm9000a_inst_avalon_slave_0_readdata,
      niosII_system_burst_16_downstream_address_to_slave => niosII_system_burst_16_downstream_address_to_slave,
      niosII_system_burst_16_downstream_arbitrationshare => niosII_system_burst_16_downstream_arbitrationshare,
      niosII_system_burst_16_downstream_burstcount => niosII_system_burst_16_downstream_burstcount,
      niosII_system_burst_16_downstream_latency_counter => niosII_system_burst_16_downstream_latency_counter,
      niosII_system_burst_16_downstream_nativeaddress => niosII_system_burst_16_downstream_nativeaddress,
      niosII_system_burst_16_downstream_read => niosII_system_burst_16_downstream_read,
      niosII_system_burst_16_downstream_write => niosII_system_burst_16_downstream_write,
      niosII_system_burst_16_downstream_writedata => niosII_system_burst_16_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_dm9000a_inst, which is an e_ptf_instance
  the_dm9000a_inst : dm9000a_inst
    port map(
      ENET_CMD => internal_ENET_CMD_from_the_dm9000a_inst,
      ENET_CS_N => internal_ENET_CS_N_from_the_dm9000a_inst,
      ENET_DATA => ENET_DATA_to_and_from_the_dm9000a_inst,
      ENET_RD_N => internal_ENET_RD_N_from_the_dm9000a_inst,
      ENET_RST_N => internal_ENET_RST_N_from_the_dm9000a_inst,
      ENET_WR_N => internal_ENET_WR_N_from_the_dm9000a_inst,
      oDATA => dm9000a_inst_avalon_slave_0_readdata,
      oINT => dm9000a_inst_avalon_slave_0_irq,
      ENET_INT => ENET_INT_to_the_dm9000a_inst,
      iCMD => dm9000a_inst_avalon_slave_0_address,
      iCS_N => dm9000a_inst_avalon_slave_0_chipselect_n,
      iDATA => dm9000a_inst_avalon_slave_0_writedata,
      iRD_N => dm9000a_inst_avalon_slave_0_read_n,
      iRST_N => dm9000a_inst_avalon_slave_0_reset_n,
      iWR_N => dm9000a_inst_avalon_slave_0_write_n
    );


  --the_high_res_timer_s1, which is an e_instance
  the_high_res_timer_s1 : high_res_timer_s1_arbitrator
    port map(
      d1_high_res_timer_s1_end_xfer => d1_high_res_timer_s1_end_xfer,
      high_res_timer_s1_address => high_res_timer_s1_address,
      high_res_timer_s1_chipselect => high_res_timer_s1_chipselect,
      high_res_timer_s1_irq_from_sa => high_res_timer_s1_irq_from_sa,
      high_res_timer_s1_readdata_from_sa => high_res_timer_s1_readdata_from_sa,
      high_res_timer_s1_reset_n => high_res_timer_s1_reset_n,
      high_res_timer_s1_write_n => high_res_timer_s1_write_n,
      high_res_timer_s1_writedata => high_res_timer_s1_writedata,
      niosII_system_burst_15_downstream_granted_high_res_timer_s1 => niosII_system_burst_15_downstream_granted_high_res_timer_s1,
      niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 => niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1,
      niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1 => niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1,
      niosII_system_burst_15_downstream_requests_high_res_timer_s1 => niosII_system_burst_15_downstream_requests_high_res_timer_s1,
      clk => internal_altpll_inst_c1_out,
      high_res_timer_s1_irq => high_res_timer_s1_irq,
      high_res_timer_s1_readdata => high_res_timer_s1_readdata,
      niosII_system_burst_15_downstream_address_to_slave => niosII_system_burst_15_downstream_address_to_slave,
      niosII_system_burst_15_downstream_arbitrationshare => niosII_system_burst_15_downstream_arbitrationshare,
      niosII_system_burst_15_downstream_burstcount => niosII_system_burst_15_downstream_burstcount,
      niosII_system_burst_15_downstream_latency_counter => niosII_system_burst_15_downstream_latency_counter,
      niosII_system_burst_15_downstream_nativeaddress => niosII_system_burst_15_downstream_nativeaddress,
      niosII_system_burst_15_downstream_read => niosII_system_burst_15_downstream_read,
      niosII_system_burst_15_downstream_write => niosII_system_burst_15_downstream_write,
      niosII_system_burst_15_downstream_writedata => niosII_system_burst_15_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_high_res_timer, which is an e_ptf_instance
  the_high_res_timer : high_res_timer
    port map(
      irq => high_res_timer_s1_irq,
      readdata => high_res_timer_s1_readdata,
      address => high_res_timer_s1_address,
      chipselect => high_res_timer_s1_chipselect,
      clk => internal_altpll_inst_c1_out,
      reset_n => high_res_timer_s1_reset_n,
      write_n => high_res_timer_s1_write_n,
      writedata => high_res_timer_s1_writedata
    );


  --the_jtag_uart_avalon_jtag_slave, which is an e_instance
  the_jtag_uart_avalon_jtag_slave : jtag_uart_avalon_jtag_slave_arbitrator
    port map(
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      jtag_uart_avalon_jtag_slave_address => jtag_uart_avalon_jtag_slave_address,
      jtag_uart_avalon_jtag_slave_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      jtag_uart_avalon_jtag_slave_dataavailable_from_sa => jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      jtag_uart_avalon_jtag_slave_read_n => jtag_uart_avalon_jtag_slave_read_n,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_readyfordata_from_sa => jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
      jtag_uart_avalon_jtag_slave_reset_n => jtag_uart_avalon_jtag_slave_reset_n,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      jtag_uart_avalon_jtag_slave_write_n => jtag_uart_avalon_jtag_slave_write_n,
      jtag_uart_avalon_jtag_slave_writedata => jtag_uart_avalon_jtag_slave_writedata,
      niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave => niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave,
      niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave => niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave,
      niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave => niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave,
      niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave => niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave,
      clk => internal_altpll_inst_c1_out,
      jtag_uart_avalon_jtag_slave_dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      jtag_uart_avalon_jtag_slave_irq => jtag_uart_avalon_jtag_slave_irq,
      jtag_uart_avalon_jtag_slave_readdata => jtag_uart_avalon_jtag_slave_readdata,
      jtag_uart_avalon_jtag_slave_readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      jtag_uart_avalon_jtag_slave_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      niosII_system_burst_6_downstream_address_to_slave => niosII_system_burst_6_downstream_address_to_slave,
      niosII_system_burst_6_downstream_arbitrationshare => niosII_system_burst_6_downstream_arbitrationshare,
      niosII_system_burst_6_downstream_burstcount => niosII_system_burst_6_downstream_burstcount,
      niosII_system_burst_6_downstream_latency_counter => niosII_system_burst_6_downstream_latency_counter,
      niosII_system_burst_6_downstream_nativeaddress => niosII_system_burst_6_downstream_nativeaddress,
      niosII_system_burst_6_downstream_read => niosII_system_burst_6_downstream_read,
      niosII_system_burst_6_downstream_write => niosII_system_burst_6_downstream_write,
      niosII_system_burst_6_downstream_writedata => niosII_system_burst_6_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_jtag_uart, which is an e_ptf_instance
  the_jtag_uart : jtag_uart
    port map(
      av_irq => jtag_uart_avalon_jtag_slave_irq,
      av_readdata => jtag_uart_avalon_jtag_slave_readdata,
      av_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      av_address => jtag_uart_avalon_jtag_slave_address,
      av_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      av_read_n => jtag_uart_avalon_jtag_slave_read_n,
      av_write_n => jtag_uart_avalon_jtag_slave_write_n,
      av_writedata => jtag_uart_avalon_jtag_slave_writedata,
      clk => internal_altpll_inst_c1_out,
      rst_n => jtag_uart_avalon_jtag_slave_reset_n
    );


  --the_lcd_display_control_slave, which is an e_instance
  the_lcd_display_control_slave : lcd_display_control_slave_arbitrator
    port map(
      d1_lcd_display_control_slave_end_xfer => d1_lcd_display_control_slave_end_xfer,
      lcd_display_control_slave_address => lcd_display_control_slave_address,
      lcd_display_control_slave_begintransfer => lcd_display_control_slave_begintransfer,
      lcd_display_control_slave_read => lcd_display_control_slave_read,
      lcd_display_control_slave_readdata_from_sa => lcd_display_control_slave_readdata_from_sa,
      lcd_display_control_slave_wait_counter_eq_0 => lcd_display_control_slave_wait_counter_eq_0,
      lcd_display_control_slave_write => lcd_display_control_slave_write,
      lcd_display_control_slave_writedata => lcd_display_control_slave_writedata,
      niosII_system_burst_7_downstream_granted_lcd_display_control_slave => niosII_system_burst_7_downstream_granted_lcd_display_control_slave,
      niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave => niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave,
      niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave => niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave,
      niosII_system_burst_7_downstream_requests_lcd_display_control_slave => niosII_system_burst_7_downstream_requests_lcd_display_control_slave,
      clk => internal_altpll_inst_c1_out,
      lcd_display_control_slave_readdata => lcd_display_control_slave_readdata,
      niosII_system_burst_7_downstream_address_to_slave => niosII_system_burst_7_downstream_address_to_slave,
      niosII_system_burst_7_downstream_arbitrationshare => niosII_system_burst_7_downstream_arbitrationshare,
      niosII_system_burst_7_downstream_burstcount => niosII_system_burst_7_downstream_burstcount,
      niosII_system_burst_7_downstream_byteenable => niosII_system_burst_7_downstream_byteenable,
      niosII_system_burst_7_downstream_latency_counter => niosII_system_burst_7_downstream_latency_counter,
      niosII_system_burst_7_downstream_nativeaddress => niosII_system_burst_7_downstream_nativeaddress,
      niosII_system_burst_7_downstream_read => niosII_system_burst_7_downstream_read,
      niosII_system_burst_7_downstream_write => niosII_system_burst_7_downstream_write,
      niosII_system_burst_7_downstream_writedata => niosII_system_burst_7_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_lcd_display, which is an e_ptf_instance
  the_lcd_display : lcd_display
    port map(
      LCD_E => internal_LCD_E_from_the_lcd_display,
      LCD_RS => internal_LCD_RS_from_the_lcd_display,
      LCD_RW => internal_LCD_RW_from_the_lcd_display,
      LCD_data => LCD_data_to_and_from_the_lcd_display,
      readdata => lcd_display_control_slave_readdata,
      address => lcd_display_control_slave_address,
      begintransfer => lcd_display_control_slave_begintransfer,
      read => lcd_display_control_slave_read,
      write => lcd_display_control_slave_write,
      writedata => lcd_display_control_slave_writedata
    );


  --the_led_pio_s1, which is an e_instance
  the_led_pio_s1 : led_pio_s1_arbitrator
    port map(
      d1_led_pio_s1_end_xfer => d1_led_pio_s1_end_xfer,
      led_pio_s1_address => led_pio_s1_address,
      led_pio_s1_chipselect => led_pio_s1_chipselect,
      led_pio_s1_readdata_from_sa => led_pio_s1_readdata_from_sa,
      led_pio_s1_reset_n => led_pio_s1_reset_n,
      led_pio_s1_write_n => led_pio_s1_write_n,
      led_pio_s1_writedata => led_pio_s1_writedata,
      niosII_system_burst_8_downstream_granted_led_pio_s1 => niosII_system_burst_8_downstream_granted_led_pio_s1,
      niosII_system_burst_8_downstream_qualified_request_led_pio_s1 => niosII_system_burst_8_downstream_qualified_request_led_pio_s1,
      niosII_system_burst_8_downstream_read_data_valid_led_pio_s1 => niosII_system_burst_8_downstream_read_data_valid_led_pio_s1,
      niosII_system_burst_8_downstream_requests_led_pio_s1 => niosII_system_burst_8_downstream_requests_led_pio_s1,
      clk => internal_altpll_inst_c1_out,
      led_pio_s1_readdata => led_pio_s1_readdata,
      niosII_system_burst_8_downstream_address_to_slave => niosII_system_burst_8_downstream_address_to_slave,
      niosII_system_burst_8_downstream_arbitrationshare => niosII_system_burst_8_downstream_arbitrationshare,
      niosII_system_burst_8_downstream_burstcount => niosII_system_burst_8_downstream_burstcount,
      niosII_system_burst_8_downstream_byteenable => niosII_system_burst_8_downstream_byteenable,
      niosII_system_burst_8_downstream_latency_counter => niosII_system_burst_8_downstream_latency_counter,
      niosII_system_burst_8_downstream_nativeaddress => niosII_system_burst_8_downstream_nativeaddress,
      niosII_system_burst_8_downstream_read => niosII_system_burst_8_downstream_read,
      niosII_system_burst_8_downstream_write => niosII_system_burst_8_downstream_write,
      niosII_system_burst_8_downstream_writedata => niosII_system_burst_8_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_led_pio, which is an e_ptf_instance
  the_led_pio : led_pio
    port map(
      out_port => internal_out_port_from_the_led_pio,
      readdata => led_pio_s1_readdata,
      address => led_pio_s1_address,
      chipselect => led_pio_s1_chipselect,
      clk => internal_altpll_inst_c1_out,
      reset_n => led_pio_s1_reset_n,
      write_n => led_pio_s1_write_n,
      writedata => led_pio_s1_writedata
    );


  --the_memory_s1, which is an e_instance
  the_memory_s1 : memory_s1_arbitrator
    port map(
      d1_memory_s1_end_xfer => d1_memory_s1_end_xfer,
      memory_s1_address => memory_s1_address,
      memory_s1_byteenable => memory_s1_byteenable,
      memory_s1_chipselect => memory_s1_chipselect,
      memory_s1_clken => memory_s1_clken,
      memory_s1_readdata_from_sa => memory_s1_readdata_from_sa,
      memory_s1_reset => memory_s1_reset,
      memory_s1_write => memory_s1_write,
      memory_s1_writedata => memory_s1_writedata,
      niosII_system_burst_2_downstream_granted_memory_s1 => niosII_system_burst_2_downstream_granted_memory_s1,
      niosII_system_burst_2_downstream_qualified_request_memory_s1 => niosII_system_burst_2_downstream_qualified_request_memory_s1,
      niosII_system_burst_2_downstream_read_data_valid_memory_s1 => niosII_system_burst_2_downstream_read_data_valid_memory_s1,
      niosII_system_burst_2_downstream_requests_memory_s1 => niosII_system_burst_2_downstream_requests_memory_s1,
      niosII_system_burst_3_downstream_granted_memory_s1 => niosII_system_burst_3_downstream_granted_memory_s1,
      niosII_system_burst_3_downstream_qualified_request_memory_s1 => niosII_system_burst_3_downstream_qualified_request_memory_s1,
      niosII_system_burst_3_downstream_read_data_valid_memory_s1 => niosII_system_burst_3_downstream_read_data_valid_memory_s1,
      niosII_system_burst_3_downstream_requests_memory_s1 => niosII_system_burst_3_downstream_requests_memory_s1,
      clk => internal_altpll_inst_c1_out,
      memory_s1_readdata => memory_s1_readdata,
      niosII_system_burst_2_downstream_address_to_slave => niosII_system_burst_2_downstream_address_to_slave,
      niosII_system_burst_2_downstream_arbitrationshare => niosII_system_burst_2_downstream_arbitrationshare,
      niosII_system_burst_2_downstream_burstcount => niosII_system_burst_2_downstream_burstcount,
      niosII_system_burst_2_downstream_byteenable => niosII_system_burst_2_downstream_byteenable,
      niosII_system_burst_2_downstream_latency_counter => niosII_system_burst_2_downstream_latency_counter,
      niosII_system_burst_2_downstream_read => niosII_system_burst_2_downstream_read,
      niosII_system_burst_2_downstream_write => niosII_system_burst_2_downstream_write,
      niosII_system_burst_2_downstream_writedata => niosII_system_burst_2_downstream_writedata,
      niosII_system_burst_3_downstream_address_to_slave => niosII_system_burst_3_downstream_address_to_slave,
      niosII_system_burst_3_downstream_arbitrationshare => niosII_system_burst_3_downstream_arbitrationshare,
      niosII_system_burst_3_downstream_burstcount => niosII_system_burst_3_downstream_burstcount,
      niosII_system_burst_3_downstream_byteenable => niosII_system_burst_3_downstream_byteenable,
      niosII_system_burst_3_downstream_latency_counter => niosII_system_burst_3_downstream_latency_counter,
      niosII_system_burst_3_downstream_read => niosII_system_burst_3_downstream_read,
      niosII_system_burst_3_downstream_write => niosII_system_burst_3_downstream_write,
      niosII_system_burst_3_downstream_writedata => niosII_system_burst_3_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_memory, which is an e_ptf_instance
  the_memory : memory
    port map(
      readdata => memory_s1_readdata,
      address => memory_s1_address,
      byteenable => memory_s1_byteenable,
      chipselect => memory_s1_chipselect,
      clk => internal_altpll_inst_c1_out,
      clken => memory_s1_clken,
      reset => memory_s1_reset,
      write => memory_s1_write,
      writedata => memory_s1_writedata
    );


  --the_niosII_system_burst_0_upstream, which is an e_instance
  the_niosII_system_burst_0_upstream : niosII_system_burst_0_upstream_arbitrator
    port map(
      cpu_instruction_master_granted_niosII_system_burst_0_upstream => cpu_instruction_master_granted_niosII_system_burst_0_upstream,
      cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream => cpu_instruction_master_qualified_request_niosII_system_burst_0_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream => cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register,
      cpu_instruction_master_requests_niosII_system_burst_0_upstream => cpu_instruction_master_requests_niosII_system_burst_0_upstream,
      d1_niosII_system_burst_0_upstream_end_xfer => d1_niosII_system_burst_0_upstream_end_xfer,
      niosII_system_burst_0_upstream_address => niosII_system_burst_0_upstream_address,
      niosII_system_burst_0_upstream_byteaddress => niosII_system_burst_0_upstream_byteaddress,
      niosII_system_burst_0_upstream_byteenable => niosII_system_burst_0_upstream_byteenable,
      niosII_system_burst_0_upstream_debugaccess => niosII_system_burst_0_upstream_debugaccess,
      niosII_system_burst_0_upstream_read => niosII_system_burst_0_upstream_read,
      niosII_system_burst_0_upstream_readdata_from_sa => niosII_system_burst_0_upstream_readdata_from_sa,
      niosII_system_burst_0_upstream_waitrequest_from_sa => niosII_system_burst_0_upstream_waitrequest_from_sa,
      niosII_system_burst_0_upstream_write => niosII_system_burst_0_upstream_write,
      clk => internal_altpll_inst_c1_out,
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_burstcount => cpu_instruction_master_burstcount,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register,
      niosII_system_burst_0_upstream_readdata => niosII_system_burst_0_upstream_readdata,
      niosII_system_burst_0_upstream_readdatavalid => niosII_system_burst_0_upstream_readdatavalid,
      niosII_system_burst_0_upstream_waitrequest => niosII_system_burst_0_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_0_downstream, which is an e_instance
  the_niosII_system_burst_0_downstream : niosII_system_burst_0_downstream_arbitrator
    port map(
      niosII_system_burst_0_downstream_address_to_slave => niosII_system_burst_0_downstream_address_to_slave,
      niosII_system_burst_0_downstream_latency_counter => niosII_system_burst_0_downstream_latency_counter,
      niosII_system_burst_0_downstream_readdata => niosII_system_burst_0_downstream_readdata,
      niosII_system_burst_0_downstream_readdatavalid => niosII_system_burst_0_downstream_readdatavalid,
      niosII_system_burst_0_downstream_reset_n => niosII_system_burst_0_downstream_reset_n,
      niosII_system_burst_0_downstream_waitrequest => niosII_system_burst_0_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      cpu_jtag_debug_module_readdata_from_sa => cpu_jtag_debug_module_readdata_from_sa,
      d1_cpu_jtag_debug_module_end_xfer => d1_cpu_jtag_debug_module_end_xfer,
      niosII_system_burst_0_downstream_address => niosII_system_burst_0_downstream_address,
      niosII_system_burst_0_downstream_burstcount => niosII_system_burst_0_downstream_burstcount,
      niosII_system_burst_0_downstream_byteenable => niosII_system_burst_0_downstream_byteenable,
      niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module => niosII_system_burst_0_downstream_granted_cpu_jtag_debug_module,
      niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module => niosII_system_burst_0_downstream_qualified_request_cpu_jtag_debug_module,
      niosII_system_burst_0_downstream_read => niosII_system_burst_0_downstream_read,
      niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module => niosII_system_burst_0_downstream_read_data_valid_cpu_jtag_debug_module,
      niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module => niosII_system_burst_0_downstream_requests_cpu_jtag_debug_module,
      niosII_system_burst_0_downstream_write => niosII_system_burst_0_downstream_write,
      niosII_system_burst_0_downstream_writedata => niosII_system_burst_0_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_0, which is an e_ptf_instance
  the_niosII_system_burst_0 : niosII_system_burst_0
    port map(
      reg_downstream_address => niosII_system_burst_0_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_0_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_0_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_0_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_0_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_0_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_0_downstream_read,
      reg_downstream_write => niosII_system_burst_0_downstream_write,
      reg_downstream_writedata => niosII_system_burst_0_downstream_writedata,
      upstream_readdata => niosII_system_burst_0_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_0_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_0_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_0_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_0_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_0_downstream_waitrequest,
      reset_n => niosII_system_burst_0_downstream_reset_n,
      upstream_address => niosII_system_burst_0_upstream_byteaddress,
      upstream_byteenable => niosII_system_burst_0_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_0_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_0_upstream_address,
      upstream_read => niosII_system_burst_0_upstream_read,
      upstream_write => niosII_system_burst_0_upstream_write,
      upstream_writedata => niosII_system_burst_0_upstream_writedata
    );


  --the_niosII_system_burst_1_upstream, which is an e_instance
  the_niosII_system_burst_1_upstream : niosII_system_burst_1_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_1_upstream => cpu_data_master_granted_niosII_system_burst_1_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_1_upstream => cpu_data_master_qualified_request_niosII_system_burst_1_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_1_upstream => cpu_data_master_requests_niosII_system_burst_1_upstream,
      d1_niosII_system_burst_1_upstream_end_xfer => d1_niosII_system_burst_1_upstream_end_xfer,
      niosII_system_burst_1_upstream_address => niosII_system_burst_1_upstream_address,
      niosII_system_burst_1_upstream_burstcount => niosII_system_burst_1_upstream_burstcount,
      niosII_system_burst_1_upstream_byteaddress => niosII_system_burst_1_upstream_byteaddress,
      niosII_system_burst_1_upstream_byteenable => niosII_system_burst_1_upstream_byteenable,
      niosII_system_burst_1_upstream_debugaccess => niosII_system_burst_1_upstream_debugaccess,
      niosII_system_burst_1_upstream_read => niosII_system_burst_1_upstream_read,
      niosII_system_burst_1_upstream_readdata_from_sa => niosII_system_burst_1_upstream_readdata_from_sa,
      niosII_system_burst_1_upstream_waitrequest_from_sa => niosII_system_burst_1_upstream_waitrequest_from_sa,
      niosII_system_burst_1_upstream_write => niosII_system_burst_1_upstream_write,
      niosII_system_burst_1_upstream_writedata => niosII_system_burst_1_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_1_upstream_readdata => niosII_system_burst_1_upstream_readdata,
      niosII_system_burst_1_upstream_readdatavalid => niosII_system_burst_1_upstream_readdatavalid,
      niosII_system_burst_1_upstream_waitrequest => niosII_system_burst_1_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_1_downstream, which is an e_instance
  the_niosII_system_burst_1_downstream : niosII_system_burst_1_downstream_arbitrator
    port map(
      niosII_system_burst_1_downstream_address_to_slave => niosII_system_burst_1_downstream_address_to_slave,
      niosII_system_burst_1_downstream_latency_counter => niosII_system_burst_1_downstream_latency_counter,
      niosII_system_burst_1_downstream_readdata => niosII_system_burst_1_downstream_readdata,
      niosII_system_burst_1_downstream_readdatavalid => niosII_system_burst_1_downstream_readdatavalid,
      niosII_system_burst_1_downstream_reset_n => niosII_system_burst_1_downstream_reset_n,
      niosII_system_burst_1_downstream_waitrequest => niosII_system_burst_1_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      cpu_jtag_debug_module_readdata_from_sa => cpu_jtag_debug_module_readdata_from_sa,
      d1_cpu_jtag_debug_module_end_xfer => d1_cpu_jtag_debug_module_end_xfer,
      niosII_system_burst_1_downstream_address => niosII_system_burst_1_downstream_address,
      niosII_system_burst_1_downstream_burstcount => niosII_system_burst_1_downstream_burstcount,
      niosII_system_burst_1_downstream_byteenable => niosII_system_burst_1_downstream_byteenable,
      niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module => niosII_system_burst_1_downstream_granted_cpu_jtag_debug_module,
      niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module => niosII_system_burst_1_downstream_qualified_request_cpu_jtag_debug_module,
      niosII_system_burst_1_downstream_read => niosII_system_burst_1_downstream_read,
      niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module => niosII_system_burst_1_downstream_read_data_valid_cpu_jtag_debug_module,
      niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module => niosII_system_burst_1_downstream_requests_cpu_jtag_debug_module,
      niosII_system_burst_1_downstream_write => niosII_system_burst_1_downstream_write,
      niosII_system_burst_1_downstream_writedata => niosII_system_burst_1_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_1, which is an e_ptf_instance
  the_niosII_system_burst_1 : niosII_system_burst_1
    port map(
      reg_downstream_address => niosII_system_burst_1_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_1_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_1_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_1_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_1_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_1_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_1_downstream_read,
      reg_downstream_write => niosII_system_burst_1_downstream_write,
      reg_downstream_writedata => niosII_system_burst_1_downstream_writedata,
      upstream_readdata => niosII_system_burst_1_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_1_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_1_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_1_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_1_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_1_downstream_waitrequest,
      reset_n => niosII_system_burst_1_downstream_reset_n,
      upstream_address => niosII_system_burst_1_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_1_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_1_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_1_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_1_upstream_address,
      upstream_read => niosII_system_burst_1_upstream_read,
      upstream_write => niosII_system_burst_1_upstream_write,
      upstream_writedata => niosII_system_burst_1_upstream_writedata
    );


  --the_niosII_system_burst_10_upstream, which is an e_instance
  the_niosII_system_burst_10_upstream : niosII_system_burst_10_upstream_arbitrator
    port map(
      cpu_instruction_master_granted_niosII_system_burst_10_upstream => cpu_instruction_master_granted_niosII_system_burst_10_upstream,
      cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream => cpu_instruction_master_qualified_request_niosII_system_burst_10_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream => cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register,
      cpu_instruction_master_requests_niosII_system_burst_10_upstream => cpu_instruction_master_requests_niosII_system_burst_10_upstream,
      d1_niosII_system_burst_10_upstream_end_xfer => d1_niosII_system_burst_10_upstream_end_xfer,
      niosII_system_burst_10_upstream_address => niosII_system_burst_10_upstream_address,
      niosII_system_burst_10_upstream_byteaddress => niosII_system_burst_10_upstream_byteaddress,
      niosII_system_burst_10_upstream_byteenable => niosII_system_burst_10_upstream_byteenable,
      niosII_system_burst_10_upstream_debugaccess => niosII_system_burst_10_upstream_debugaccess,
      niosII_system_burst_10_upstream_read => niosII_system_burst_10_upstream_read,
      niosII_system_burst_10_upstream_readdata_from_sa => niosII_system_burst_10_upstream_readdata_from_sa,
      niosII_system_burst_10_upstream_waitrequest_from_sa => niosII_system_burst_10_upstream_waitrequest_from_sa,
      niosII_system_burst_10_upstream_write => niosII_system_burst_10_upstream_write,
      clk => internal_altpll_inst_c1_out,
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_burstcount => cpu_instruction_master_burstcount,
      cpu_instruction_master_dbs_address => cpu_instruction_master_dbs_address,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register,
      niosII_system_burst_10_upstream_readdata => niosII_system_burst_10_upstream_readdata,
      niosII_system_burst_10_upstream_readdatavalid => niosII_system_burst_10_upstream_readdatavalid,
      niosII_system_burst_10_upstream_waitrequest => niosII_system_burst_10_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_10_downstream, which is an e_instance
  the_niosII_system_burst_10_downstream : niosII_system_burst_10_downstream_arbitrator
    port map(
      niosII_system_burst_10_downstream_address_to_slave => niosII_system_burst_10_downstream_address_to_slave,
      niosII_system_burst_10_downstream_latency_counter => niosII_system_burst_10_downstream_latency_counter,
      niosII_system_burst_10_downstream_readdata => niosII_system_burst_10_downstream_readdata,
      niosII_system_burst_10_downstream_readdatavalid => niosII_system_burst_10_downstream_readdatavalid,
      niosII_system_burst_10_downstream_reset_n => niosII_system_burst_10_downstream_reset_n,
      niosII_system_burst_10_downstream_waitrequest => niosII_system_burst_10_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      niosII_system_burst_10_downstream_address => niosII_system_burst_10_downstream_address,
      niosII_system_burst_10_downstream_burstcount => niosII_system_burst_10_downstream_burstcount,
      niosII_system_burst_10_downstream_byteenable => niosII_system_burst_10_downstream_byteenable,
      niosII_system_burst_10_downstream_granted_sdram_s1 => niosII_system_burst_10_downstream_granted_sdram_s1,
      niosII_system_burst_10_downstream_qualified_request_sdram_s1 => niosII_system_burst_10_downstream_qualified_request_sdram_s1,
      niosII_system_burst_10_downstream_read => niosII_system_burst_10_downstream_read,
      niosII_system_burst_10_downstream_read_data_valid_sdram_s1 => niosII_system_burst_10_downstream_read_data_valid_sdram_s1,
      niosII_system_burst_10_downstream_read_data_valid_sdram_s1_shift_register => niosII_system_burst_10_downstream_read_data_valid_sdram_s1_shift_register,
      niosII_system_burst_10_downstream_requests_sdram_s1 => niosII_system_burst_10_downstream_requests_sdram_s1,
      niosII_system_burst_10_downstream_write => niosII_system_burst_10_downstream_write,
      niosII_system_burst_10_downstream_writedata => niosII_system_burst_10_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa
    );


  --the_niosII_system_burst_10, which is an e_ptf_instance
  the_niosII_system_burst_10 : niosII_system_burst_10
    port map(
      reg_downstream_address => niosII_system_burst_10_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_10_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_10_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_10_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_10_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_10_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_10_downstream_read,
      reg_downstream_write => niosII_system_burst_10_downstream_write,
      reg_downstream_writedata => niosII_system_burst_10_downstream_writedata,
      upstream_readdata => niosII_system_burst_10_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_10_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_10_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_10_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_10_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_10_downstream_waitrequest,
      reset_n => niosII_system_burst_10_downstream_reset_n,
      upstream_address => niosII_system_burst_10_upstream_byteaddress,
      upstream_byteenable => niosII_system_burst_10_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_10_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_10_upstream_address,
      upstream_read => niosII_system_burst_10_upstream_read,
      upstream_write => niosII_system_burst_10_upstream_write,
      upstream_writedata => niosII_system_burst_10_upstream_writedata
    );


  --the_niosII_system_burst_11_upstream, which is an e_instance
  the_niosII_system_burst_11_upstream : niosII_system_burst_11_upstream_arbitrator
    port map(
      cpu_data_master_byteenable_niosII_system_burst_11_upstream => cpu_data_master_byteenable_niosII_system_burst_11_upstream,
      cpu_data_master_granted_niosII_system_burst_11_upstream => cpu_data_master_granted_niosII_system_burst_11_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_11_upstream => cpu_data_master_qualified_request_niosII_system_burst_11_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_11_upstream => cpu_data_master_requests_niosII_system_burst_11_upstream,
      d1_niosII_system_burst_11_upstream_end_xfer => d1_niosII_system_burst_11_upstream_end_xfer,
      niosII_system_burst_11_upstream_address => niosII_system_burst_11_upstream_address,
      niosII_system_burst_11_upstream_burstcount => niosII_system_burst_11_upstream_burstcount,
      niosII_system_burst_11_upstream_byteaddress => niosII_system_burst_11_upstream_byteaddress,
      niosII_system_burst_11_upstream_byteenable => niosII_system_burst_11_upstream_byteenable,
      niosII_system_burst_11_upstream_debugaccess => niosII_system_burst_11_upstream_debugaccess,
      niosII_system_burst_11_upstream_read => niosII_system_burst_11_upstream_read,
      niosII_system_burst_11_upstream_readdata_from_sa => niosII_system_burst_11_upstream_readdata_from_sa,
      niosII_system_burst_11_upstream_waitrequest_from_sa => niosII_system_burst_11_upstream_waitrequest_from_sa,
      niosII_system_burst_11_upstream_write => niosII_system_burst_11_upstream_write,
      niosII_system_burst_11_upstream_writedata => niosII_system_burst_11_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_dbs_address => cpu_data_master_dbs_address,
      cpu_data_master_dbs_write_16 => cpu_data_master_dbs_write_16,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      niosII_system_burst_11_upstream_readdata => niosII_system_burst_11_upstream_readdata,
      niosII_system_burst_11_upstream_readdatavalid => niosII_system_burst_11_upstream_readdatavalid,
      niosII_system_burst_11_upstream_waitrequest => niosII_system_burst_11_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_11_downstream, which is an e_instance
  the_niosII_system_burst_11_downstream : niosII_system_burst_11_downstream_arbitrator
    port map(
      niosII_system_burst_11_downstream_address_to_slave => niosII_system_burst_11_downstream_address_to_slave,
      niosII_system_burst_11_downstream_latency_counter => niosII_system_burst_11_downstream_latency_counter,
      niosII_system_burst_11_downstream_readdata => niosII_system_burst_11_downstream_readdata,
      niosII_system_burst_11_downstream_readdatavalid => niosII_system_burst_11_downstream_readdatavalid,
      niosII_system_burst_11_downstream_reset_n => niosII_system_burst_11_downstream_reset_n,
      niosII_system_burst_11_downstream_waitrequest => niosII_system_burst_11_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      niosII_system_burst_11_downstream_address => niosII_system_burst_11_downstream_address,
      niosII_system_burst_11_downstream_burstcount => niosII_system_burst_11_downstream_burstcount,
      niosII_system_burst_11_downstream_byteenable => niosII_system_burst_11_downstream_byteenable,
      niosII_system_burst_11_downstream_granted_sdram_s1 => niosII_system_burst_11_downstream_granted_sdram_s1,
      niosII_system_burst_11_downstream_qualified_request_sdram_s1 => niosII_system_burst_11_downstream_qualified_request_sdram_s1,
      niosII_system_burst_11_downstream_read => niosII_system_burst_11_downstream_read,
      niosII_system_burst_11_downstream_read_data_valid_sdram_s1 => niosII_system_burst_11_downstream_read_data_valid_sdram_s1,
      niosII_system_burst_11_downstream_read_data_valid_sdram_s1_shift_register => niosII_system_burst_11_downstream_read_data_valid_sdram_s1_shift_register,
      niosII_system_burst_11_downstream_requests_sdram_s1 => niosII_system_burst_11_downstream_requests_sdram_s1,
      niosII_system_burst_11_downstream_write => niosII_system_burst_11_downstream_write,
      niosII_system_burst_11_downstream_writedata => niosII_system_burst_11_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa
    );


  --the_niosII_system_burst_11, which is an e_ptf_instance
  the_niosII_system_burst_11 : niosII_system_burst_11
    port map(
      reg_downstream_address => niosII_system_burst_11_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_11_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_11_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_11_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_11_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_11_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_11_downstream_read,
      reg_downstream_write => niosII_system_burst_11_downstream_write,
      reg_downstream_writedata => niosII_system_burst_11_downstream_writedata,
      upstream_readdata => niosII_system_burst_11_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_11_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_11_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_11_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_11_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_11_downstream_waitrequest,
      reset_n => niosII_system_burst_11_downstream_reset_n,
      upstream_address => niosII_system_burst_11_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_11_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_11_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_11_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_11_upstream_address,
      upstream_read => niosII_system_burst_11_upstream_read,
      upstream_write => niosII_system_burst_11_upstream_write,
      upstream_writedata => niosII_system_burst_11_upstream_writedata
    );


  --the_niosII_system_burst_12_upstream, which is an e_instance
  the_niosII_system_burst_12_upstream : niosII_system_burst_12_upstream_arbitrator
    port map(
      cpu_instruction_master_granted_niosII_system_burst_12_upstream => cpu_instruction_master_granted_niosII_system_burst_12_upstream,
      cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream => cpu_instruction_master_qualified_request_niosII_system_burst_12_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream => cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register,
      cpu_instruction_master_requests_niosII_system_burst_12_upstream => cpu_instruction_master_requests_niosII_system_burst_12_upstream,
      d1_niosII_system_burst_12_upstream_end_xfer => d1_niosII_system_burst_12_upstream_end_xfer,
      niosII_system_burst_12_upstream_address => niosII_system_burst_12_upstream_address,
      niosII_system_burst_12_upstream_byteaddress => niosII_system_burst_12_upstream_byteaddress,
      niosII_system_burst_12_upstream_byteenable => niosII_system_burst_12_upstream_byteenable,
      niosII_system_burst_12_upstream_debugaccess => niosII_system_burst_12_upstream_debugaccess,
      niosII_system_burst_12_upstream_read => niosII_system_burst_12_upstream_read,
      niosII_system_burst_12_upstream_readdata_from_sa => niosII_system_burst_12_upstream_readdata_from_sa,
      niosII_system_burst_12_upstream_waitrequest_from_sa => niosII_system_burst_12_upstream_waitrequest_from_sa,
      niosII_system_burst_12_upstream_write => niosII_system_burst_12_upstream_write,
      clk => internal_altpll_inst_c1_out,
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_burstcount => cpu_instruction_master_burstcount,
      cpu_instruction_master_dbs_address => cpu_instruction_master_dbs_address,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register,
      niosII_system_burst_12_upstream_readdata => niosII_system_burst_12_upstream_readdata,
      niosII_system_burst_12_upstream_readdatavalid => niosII_system_burst_12_upstream_readdatavalid,
      niosII_system_burst_12_upstream_waitrequest => niosII_system_burst_12_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_12_downstream, which is an e_instance
  the_niosII_system_burst_12_downstream : niosII_system_burst_12_downstream_arbitrator
    port map(
      niosII_system_burst_12_downstream_address_to_slave => niosII_system_burst_12_downstream_address_to_slave,
      niosII_system_burst_12_downstream_latency_counter => niosII_system_burst_12_downstream_latency_counter,
      niosII_system_burst_12_downstream_readdata => niosII_system_burst_12_downstream_readdata,
      niosII_system_burst_12_downstream_readdatavalid => niosII_system_burst_12_downstream_readdatavalid,
      niosII_system_burst_12_downstream_reset_n => niosII_system_burst_12_downstream_reset_n,
      niosII_system_burst_12_downstream_waitrequest => niosII_system_burst_12_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_tri_state_bridge_avalon_slave_end_xfer => d1_tri_state_bridge_avalon_slave_end_xfer,
      ext_flash_s1_wait_counter_eq_0 => ext_flash_s1_wait_counter_eq_0,
      incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 => incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0,
      niosII_system_burst_12_downstream_address => niosII_system_burst_12_downstream_address,
      niosII_system_burst_12_downstream_burstcount => niosII_system_burst_12_downstream_burstcount,
      niosII_system_burst_12_downstream_byteenable => niosII_system_burst_12_downstream_byteenable,
      niosII_system_burst_12_downstream_granted_ext_flash_s1 => niosII_system_burst_12_downstream_granted_ext_flash_s1,
      niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 => niosII_system_burst_12_downstream_qualified_request_ext_flash_s1,
      niosII_system_burst_12_downstream_read => niosII_system_burst_12_downstream_read,
      niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1 => niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1,
      niosII_system_burst_12_downstream_requests_ext_flash_s1 => niosII_system_burst_12_downstream_requests_ext_flash_s1,
      niosII_system_burst_12_downstream_write => niosII_system_burst_12_downstream_write,
      niosII_system_burst_12_downstream_writedata => niosII_system_burst_12_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_12, which is an e_ptf_instance
  the_niosII_system_burst_12 : niosII_system_burst_12
    port map(
      reg_downstream_address => niosII_system_burst_12_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_12_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_12_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_12_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_12_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_12_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_12_downstream_read,
      reg_downstream_write => niosII_system_burst_12_downstream_write,
      reg_downstream_writedata => niosII_system_burst_12_downstream_writedata,
      upstream_readdata => niosII_system_burst_12_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_12_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_12_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_12_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_12_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_12_downstream_waitrequest,
      reset_n => niosII_system_burst_12_downstream_reset_n,
      upstream_address => niosII_system_burst_12_upstream_byteaddress,
      upstream_byteenable => niosII_system_burst_12_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_12_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_12_upstream_address,
      upstream_read => niosII_system_burst_12_upstream_read,
      upstream_write => niosII_system_burst_12_upstream_write,
      upstream_writedata => niosII_system_burst_12_upstream_writedata
    );


  --the_niosII_system_burst_13_upstream, which is an e_instance
  the_niosII_system_burst_13_upstream : niosII_system_burst_13_upstream_arbitrator
    port map(
      cpu_data_master_byteenable_niosII_system_burst_13_upstream => cpu_data_master_byteenable_niosII_system_burst_13_upstream,
      cpu_data_master_granted_niosII_system_burst_13_upstream => cpu_data_master_granted_niosII_system_burst_13_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_13_upstream => cpu_data_master_qualified_request_niosII_system_burst_13_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_13_upstream => cpu_data_master_requests_niosII_system_burst_13_upstream,
      d1_niosII_system_burst_13_upstream_end_xfer => d1_niosII_system_burst_13_upstream_end_xfer,
      niosII_system_burst_13_upstream_address => niosII_system_burst_13_upstream_address,
      niosII_system_burst_13_upstream_burstcount => niosII_system_burst_13_upstream_burstcount,
      niosII_system_burst_13_upstream_byteaddress => niosII_system_burst_13_upstream_byteaddress,
      niosII_system_burst_13_upstream_byteenable => niosII_system_burst_13_upstream_byteenable,
      niosII_system_burst_13_upstream_debugaccess => niosII_system_burst_13_upstream_debugaccess,
      niosII_system_burst_13_upstream_read => niosII_system_burst_13_upstream_read,
      niosII_system_burst_13_upstream_readdata_from_sa => niosII_system_burst_13_upstream_readdata_from_sa,
      niosII_system_burst_13_upstream_waitrequest_from_sa => niosII_system_burst_13_upstream_waitrequest_from_sa,
      niosII_system_burst_13_upstream_write => niosII_system_burst_13_upstream_write,
      niosII_system_burst_13_upstream_writedata => niosII_system_burst_13_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_dbs_address => cpu_data_master_dbs_address,
      cpu_data_master_dbs_write_8 => cpu_data_master_dbs_write_8,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      niosII_system_burst_13_upstream_readdata => niosII_system_burst_13_upstream_readdata,
      niosII_system_burst_13_upstream_readdatavalid => niosII_system_burst_13_upstream_readdatavalid,
      niosII_system_burst_13_upstream_waitrequest => niosII_system_burst_13_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_13_downstream, which is an e_instance
  the_niosII_system_burst_13_downstream : niosII_system_burst_13_downstream_arbitrator
    port map(
      niosII_system_burst_13_downstream_address_to_slave => niosII_system_burst_13_downstream_address_to_slave,
      niosII_system_burst_13_downstream_latency_counter => niosII_system_burst_13_downstream_latency_counter,
      niosII_system_burst_13_downstream_readdata => niosII_system_burst_13_downstream_readdata,
      niosII_system_burst_13_downstream_readdatavalid => niosII_system_burst_13_downstream_readdatavalid,
      niosII_system_burst_13_downstream_reset_n => niosII_system_burst_13_downstream_reset_n,
      niosII_system_burst_13_downstream_waitrequest => niosII_system_burst_13_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_tri_state_bridge_avalon_slave_end_xfer => d1_tri_state_bridge_avalon_slave_end_xfer,
      ext_flash_s1_wait_counter_eq_0 => ext_flash_s1_wait_counter_eq_0,
      incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 => incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0,
      niosII_system_burst_13_downstream_address => niosII_system_burst_13_downstream_address,
      niosII_system_burst_13_downstream_burstcount => niosII_system_burst_13_downstream_burstcount,
      niosII_system_burst_13_downstream_byteenable => niosII_system_burst_13_downstream_byteenable,
      niosII_system_burst_13_downstream_granted_ext_flash_s1 => niosII_system_burst_13_downstream_granted_ext_flash_s1,
      niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 => niosII_system_burst_13_downstream_qualified_request_ext_flash_s1,
      niosII_system_burst_13_downstream_read => niosII_system_burst_13_downstream_read,
      niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1 => niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1,
      niosII_system_burst_13_downstream_requests_ext_flash_s1 => niosII_system_burst_13_downstream_requests_ext_flash_s1,
      niosII_system_burst_13_downstream_write => niosII_system_burst_13_downstream_write,
      niosII_system_burst_13_downstream_writedata => niosII_system_burst_13_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_13, which is an e_ptf_instance
  the_niosII_system_burst_13 : niosII_system_burst_13
    port map(
      reg_downstream_address => niosII_system_burst_13_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_13_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_13_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_13_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_13_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_13_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_13_downstream_read,
      reg_downstream_write => niosII_system_burst_13_downstream_write,
      reg_downstream_writedata => niosII_system_burst_13_downstream_writedata,
      upstream_readdata => niosII_system_burst_13_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_13_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_13_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_13_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_13_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_13_downstream_waitrequest,
      reset_n => niosII_system_burst_13_downstream_reset_n,
      upstream_address => niosII_system_burst_13_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_13_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_13_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_13_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_13_upstream_address,
      upstream_read => niosII_system_burst_13_upstream_read,
      upstream_write => niosII_system_burst_13_upstream_write,
      upstream_writedata => niosII_system_burst_13_upstream_writedata
    );


  --the_niosII_system_burst_14_upstream, which is an e_instance
  the_niosII_system_burst_14_upstream : niosII_system_burst_14_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_14_upstream => cpu_data_master_granted_niosII_system_burst_14_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_14_upstream => cpu_data_master_qualified_request_niosII_system_burst_14_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_14_upstream => cpu_data_master_requests_niosII_system_burst_14_upstream,
      d1_niosII_system_burst_14_upstream_end_xfer => d1_niosII_system_burst_14_upstream_end_xfer,
      niosII_system_burst_14_upstream_address => niosII_system_burst_14_upstream_address,
      niosII_system_burst_14_upstream_burstcount => niosII_system_burst_14_upstream_burstcount,
      niosII_system_burst_14_upstream_byteaddress => niosII_system_burst_14_upstream_byteaddress,
      niosII_system_burst_14_upstream_byteenable => niosII_system_burst_14_upstream_byteenable,
      niosII_system_burst_14_upstream_debugaccess => niosII_system_burst_14_upstream_debugaccess,
      niosII_system_burst_14_upstream_read => niosII_system_burst_14_upstream_read,
      niosII_system_burst_14_upstream_readdata_from_sa => niosII_system_burst_14_upstream_readdata_from_sa,
      niosII_system_burst_14_upstream_waitrequest_from_sa => niosII_system_burst_14_upstream_waitrequest_from_sa,
      niosII_system_burst_14_upstream_write => niosII_system_burst_14_upstream_write,
      niosII_system_burst_14_upstream_writedata => niosII_system_burst_14_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_14_upstream_readdata => niosII_system_burst_14_upstream_readdata,
      niosII_system_burst_14_upstream_readdatavalid => niosII_system_burst_14_upstream_readdatavalid,
      niosII_system_burst_14_upstream_waitrequest => niosII_system_burst_14_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_14_downstream, which is an e_instance
  the_niosII_system_burst_14_downstream : niosII_system_burst_14_downstream_arbitrator
    port map(
      niosII_system_burst_14_downstream_address_to_slave => niosII_system_burst_14_downstream_address_to_slave,
      niosII_system_burst_14_downstream_latency_counter => niosII_system_burst_14_downstream_latency_counter,
      niosII_system_burst_14_downstream_readdata => niosII_system_burst_14_downstream_readdata,
      niosII_system_burst_14_downstream_readdatavalid => niosII_system_burst_14_downstream_readdatavalid,
      niosII_system_burst_14_downstream_reset_n => niosII_system_burst_14_downstream_reset_n,
      niosII_system_burst_14_downstream_waitrequest => niosII_system_burst_14_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_seven_seg_pio_s1_end_xfer => d1_seven_seg_pio_s1_end_xfer,
      niosII_system_burst_14_downstream_address => niosII_system_burst_14_downstream_address,
      niosII_system_burst_14_downstream_burstcount => niosII_system_burst_14_downstream_burstcount,
      niosII_system_burst_14_downstream_byteenable => niosII_system_burst_14_downstream_byteenable,
      niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 => niosII_system_burst_14_downstream_granted_seven_seg_pio_s1,
      niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 => niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1,
      niosII_system_burst_14_downstream_read => niosII_system_burst_14_downstream_read,
      niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1 => niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1,
      niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 => niosII_system_burst_14_downstream_requests_seven_seg_pio_s1,
      niosII_system_burst_14_downstream_write => niosII_system_burst_14_downstream_write,
      niosII_system_burst_14_downstream_writedata => niosII_system_burst_14_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      seven_seg_pio_s1_readdata_from_sa => seven_seg_pio_s1_readdata_from_sa
    );


  --the_niosII_system_burst_14, which is an e_ptf_instance
  the_niosII_system_burst_14 : niosII_system_burst_14
    port map(
      reg_downstream_address => niosII_system_burst_14_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_14_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_14_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_14_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_14_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_14_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_14_downstream_read,
      reg_downstream_write => niosII_system_burst_14_downstream_write,
      reg_downstream_writedata => niosII_system_burst_14_downstream_writedata,
      upstream_readdata => niosII_system_burst_14_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_14_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_14_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_14_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_14_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_14_downstream_waitrequest,
      reset_n => niosII_system_burst_14_downstream_reset_n,
      upstream_address => niosII_system_burst_14_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_14_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_14_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_14_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_14_upstream_address,
      upstream_read => niosII_system_burst_14_upstream_read,
      upstream_write => niosII_system_burst_14_upstream_write,
      upstream_writedata => niosII_system_burst_14_upstream_writedata
    );


  --the_niosII_system_burst_15_upstream, which is an e_instance
  the_niosII_system_burst_15_upstream : niosII_system_burst_15_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_15_upstream => cpu_data_master_granted_niosII_system_burst_15_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_15_upstream => cpu_data_master_qualified_request_niosII_system_burst_15_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_15_upstream => cpu_data_master_requests_niosII_system_burst_15_upstream,
      d1_niosII_system_burst_15_upstream_end_xfer => d1_niosII_system_burst_15_upstream_end_xfer,
      niosII_system_burst_15_upstream_address => niosII_system_burst_15_upstream_address,
      niosII_system_burst_15_upstream_burstcount => niosII_system_burst_15_upstream_burstcount,
      niosII_system_burst_15_upstream_byteaddress => niosII_system_burst_15_upstream_byteaddress,
      niosII_system_burst_15_upstream_byteenable => niosII_system_burst_15_upstream_byteenable,
      niosII_system_burst_15_upstream_debugaccess => niosII_system_burst_15_upstream_debugaccess,
      niosII_system_burst_15_upstream_read => niosII_system_burst_15_upstream_read,
      niosII_system_burst_15_upstream_readdata_from_sa => niosII_system_burst_15_upstream_readdata_from_sa,
      niosII_system_burst_15_upstream_waitrequest_from_sa => niosII_system_burst_15_upstream_waitrequest_from_sa,
      niosII_system_burst_15_upstream_write => niosII_system_burst_15_upstream_write,
      niosII_system_burst_15_upstream_writedata => niosII_system_burst_15_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_15_upstream_readdata => niosII_system_burst_15_upstream_readdata,
      niosII_system_burst_15_upstream_readdatavalid => niosII_system_burst_15_upstream_readdatavalid,
      niosII_system_burst_15_upstream_waitrequest => niosII_system_burst_15_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_15_downstream, which is an e_instance
  the_niosII_system_burst_15_downstream : niosII_system_burst_15_downstream_arbitrator
    port map(
      niosII_system_burst_15_downstream_address_to_slave => niosII_system_burst_15_downstream_address_to_slave,
      niosII_system_burst_15_downstream_latency_counter => niosII_system_burst_15_downstream_latency_counter,
      niosII_system_burst_15_downstream_readdata => niosII_system_burst_15_downstream_readdata,
      niosII_system_burst_15_downstream_readdatavalid => niosII_system_burst_15_downstream_readdatavalid,
      niosII_system_burst_15_downstream_reset_n => niosII_system_burst_15_downstream_reset_n,
      niosII_system_burst_15_downstream_waitrequest => niosII_system_burst_15_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_high_res_timer_s1_end_xfer => d1_high_res_timer_s1_end_xfer,
      high_res_timer_s1_readdata_from_sa => high_res_timer_s1_readdata_from_sa,
      niosII_system_burst_15_downstream_address => niosII_system_burst_15_downstream_address,
      niosII_system_burst_15_downstream_burstcount => niosII_system_burst_15_downstream_burstcount,
      niosII_system_burst_15_downstream_byteenable => niosII_system_burst_15_downstream_byteenable,
      niosII_system_burst_15_downstream_granted_high_res_timer_s1 => niosII_system_burst_15_downstream_granted_high_res_timer_s1,
      niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1 => niosII_system_burst_15_downstream_qualified_request_high_res_timer_s1,
      niosII_system_burst_15_downstream_read => niosII_system_burst_15_downstream_read,
      niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1 => niosII_system_burst_15_downstream_read_data_valid_high_res_timer_s1,
      niosII_system_burst_15_downstream_requests_high_res_timer_s1 => niosII_system_burst_15_downstream_requests_high_res_timer_s1,
      niosII_system_burst_15_downstream_write => niosII_system_burst_15_downstream_write,
      niosII_system_burst_15_downstream_writedata => niosII_system_burst_15_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_15, which is an e_ptf_instance
  the_niosII_system_burst_15 : niosII_system_burst_15
    port map(
      reg_downstream_address => niosII_system_burst_15_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_15_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_15_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_15_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_15_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_15_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_15_downstream_read,
      reg_downstream_write => niosII_system_burst_15_downstream_write,
      reg_downstream_writedata => niosII_system_burst_15_downstream_writedata,
      upstream_readdata => niosII_system_burst_15_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_15_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_15_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_15_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_15_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_15_downstream_waitrequest,
      reset_n => niosII_system_burst_15_downstream_reset_n,
      upstream_address => niosII_system_burst_15_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_15_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_15_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_15_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_15_upstream_address,
      upstream_read => niosII_system_burst_15_upstream_read,
      upstream_write => niosII_system_burst_15_upstream_write,
      upstream_writedata => niosII_system_burst_15_upstream_writedata
    );


  --the_niosII_system_burst_16_upstream, which is an e_instance
  the_niosII_system_burst_16_upstream : niosII_system_burst_16_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_16_upstream => cpu_data_master_granted_niosII_system_burst_16_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_16_upstream => cpu_data_master_qualified_request_niosII_system_burst_16_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_16_upstream => cpu_data_master_requests_niosII_system_burst_16_upstream,
      d1_niosII_system_burst_16_upstream_end_xfer => d1_niosII_system_burst_16_upstream_end_xfer,
      niosII_system_burst_16_upstream_address => niosII_system_burst_16_upstream_address,
      niosII_system_burst_16_upstream_burstcount => niosII_system_burst_16_upstream_burstcount,
      niosII_system_burst_16_upstream_byteaddress => niosII_system_burst_16_upstream_byteaddress,
      niosII_system_burst_16_upstream_byteenable => niosII_system_burst_16_upstream_byteenable,
      niosII_system_burst_16_upstream_debugaccess => niosII_system_burst_16_upstream_debugaccess,
      niosII_system_burst_16_upstream_read => niosII_system_burst_16_upstream_read,
      niosII_system_burst_16_upstream_readdata_from_sa => niosII_system_burst_16_upstream_readdata_from_sa,
      niosII_system_burst_16_upstream_waitrequest_from_sa => niosII_system_burst_16_upstream_waitrequest_from_sa,
      niosII_system_burst_16_upstream_write => niosII_system_burst_16_upstream_write,
      niosII_system_burst_16_upstream_writedata => niosII_system_burst_16_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_16_upstream_readdata => niosII_system_burst_16_upstream_readdata,
      niosII_system_burst_16_upstream_readdatavalid => niosII_system_burst_16_upstream_readdatavalid,
      niosII_system_burst_16_upstream_waitrequest => niosII_system_burst_16_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_16_downstream, which is an e_instance
  the_niosII_system_burst_16_downstream : niosII_system_burst_16_downstream_arbitrator
    port map(
      niosII_system_burst_16_downstream_address_to_slave => niosII_system_burst_16_downstream_address_to_slave,
      niosII_system_burst_16_downstream_latency_counter => niosII_system_burst_16_downstream_latency_counter,
      niosII_system_burst_16_downstream_readdata => niosII_system_burst_16_downstream_readdata,
      niosII_system_burst_16_downstream_readdatavalid => niosII_system_burst_16_downstream_readdatavalid,
      niosII_system_burst_16_downstream_reset_n => niosII_system_burst_16_downstream_reset_n,
      niosII_system_burst_16_downstream_waitrequest => niosII_system_burst_16_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_dm9000a_inst_avalon_slave_0_end_xfer => d1_dm9000a_inst_avalon_slave_0_end_xfer,
      dm9000a_inst_avalon_slave_0_readdata_from_sa => dm9000a_inst_avalon_slave_0_readdata_from_sa,
      niosII_system_burst_16_downstream_address => niosII_system_burst_16_downstream_address,
      niosII_system_burst_16_downstream_burstcount => niosII_system_burst_16_downstream_burstcount,
      niosII_system_burst_16_downstream_byteenable => niosII_system_burst_16_downstream_byteenable,
      niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0 => niosII_system_burst_16_downstream_granted_dm9000a_inst_avalon_slave_0,
      niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0 => niosII_system_burst_16_downstream_qualified_request_dm9000a_inst_avalon_slave_0,
      niosII_system_burst_16_downstream_read => niosII_system_burst_16_downstream_read,
      niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0 => niosII_system_burst_16_downstream_read_data_valid_dm9000a_inst_avalon_slave_0,
      niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0 => niosII_system_burst_16_downstream_requests_dm9000a_inst_avalon_slave_0,
      niosII_system_burst_16_downstream_write => niosII_system_burst_16_downstream_write,
      niosII_system_burst_16_downstream_writedata => niosII_system_burst_16_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_16, which is an e_ptf_instance
  the_niosII_system_burst_16 : niosII_system_burst_16
    port map(
      reg_downstream_address => niosII_system_burst_16_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_16_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_16_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_16_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_16_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_16_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_16_downstream_read,
      reg_downstream_write => niosII_system_burst_16_downstream_write,
      reg_downstream_writedata => niosII_system_burst_16_downstream_writedata,
      upstream_readdata => niosII_system_burst_16_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_16_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_16_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_16_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_16_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_16_downstream_waitrequest,
      reset_n => niosII_system_burst_16_downstream_reset_n,
      upstream_address => niosII_system_burst_16_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_16_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_16_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_16_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_16_upstream_address,
      upstream_read => niosII_system_burst_16_upstream_read,
      upstream_write => niosII_system_burst_16_upstream_write,
      upstream_writedata => niosII_system_burst_16_upstream_writedata
    );


  --the_niosII_system_burst_17_upstream, which is an e_instance
  the_niosII_system_burst_17_upstream : niosII_system_burst_17_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_17_upstream => cpu_data_master_granted_niosII_system_burst_17_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_17_upstream => cpu_data_master_qualified_request_niosII_system_burst_17_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_17_upstream => cpu_data_master_requests_niosII_system_burst_17_upstream,
      d1_niosII_system_burst_17_upstream_end_xfer => d1_niosII_system_burst_17_upstream_end_xfer,
      niosII_system_burst_17_upstream_address => niosII_system_burst_17_upstream_address,
      niosII_system_burst_17_upstream_burstcount => niosII_system_burst_17_upstream_burstcount,
      niosII_system_burst_17_upstream_byteaddress => niosII_system_burst_17_upstream_byteaddress,
      niosII_system_burst_17_upstream_byteenable => niosII_system_burst_17_upstream_byteenable,
      niosII_system_burst_17_upstream_debugaccess => niosII_system_burst_17_upstream_debugaccess,
      niosII_system_burst_17_upstream_read => niosII_system_burst_17_upstream_read,
      niosII_system_burst_17_upstream_readdata_from_sa => niosII_system_burst_17_upstream_readdata_from_sa,
      niosII_system_burst_17_upstream_waitrequest_from_sa => niosII_system_burst_17_upstream_waitrequest_from_sa,
      niosII_system_burst_17_upstream_write => niosII_system_burst_17_upstream_write,
      niosII_system_burst_17_upstream_writedata => niosII_system_burst_17_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_17_upstream_readdata => niosII_system_burst_17_upstream_readdata,
      niosII_system_burst_17_upstream_readdatavalid => niosII_system_burst_17_upstream_readdatavalid,
      niosII_system_burst_17_upstream_waitrequest => niosII_system_burst_17_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_17_downstream, which is an e_instance
  the_niosII_system_burst_17_downstream : niosII_system_burst_17_downstream_arbitrator
    port map(
      niosII_system_burst_17_downstream_address_to_slave => niosII_system_burst_17_downstream_address_to_slave,
      niosII_system_burst_17_downstream_latency_counter => niosII_system_burst_17_downstream_latency_counter,
      niosII_system_burst_17_downstream_readdata => niosII_system_burst_17_downstream_readdata,
      niosII_system_burst_17_downstream_readdatavalid => niosII_system_burst_17_downstream_readdatavalid,
      niosII_system_burst_17_downstream_reset_n => niosII_system_burst_17_downstream_reset_n,
      niosII_system_burst_17_downstream_waitrequest => niosII_system_burst_17_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_uart_0_s1_end_xfer => d1_uart_0_s1_end_xfer,
      niosII_system_burst_17_downstream_address => niosII_system_burst_17_downstream_address,
      niosII_system_burst_17_downstream_burstcount => niosII_system_burst_17_downstream_burstcount,
      niosII_system_burst_17_downstream_byteenable => niosII_system_burst_17_downstream_byteenable,
      niosII_system_burst_17_downstream_granted_uart_0_s1 => niosII_system_burst_17_downstream_granted_uart_0_s1,
      niosII_system_burst_17_downstream_qualified_request_uart_0_s1 => niosII_system_burst_17_downstream_qualified_request_uart_0_s1,
      niosII_system_burst_17_downstream_read => niosII_system_burst_17_downstream_read,
      niosII_system_burst_17_downstream_read_data_valid_uart_0_s1 => niosII_system_burst_17_downstream_read_data_valid_uart_0_s1,
      niosII_system_burst_17_downstream_requests_uart_0_s1 => niosII_system_burst_17_downstream_requests_uart_0_s1,
      niosII_system_burst_17_downstream_write => niosII_system_burst_17_downstream_write,
      niosII_system_burst_17_downstream_writedata => niosII_system_burst_17_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      uart_0_s1_readdata_from_sa => uart_0_s1_readdata_from_sa
    );


  --the_niosII_system_burst_17, which is an e_ptf_instance
  the_niosII_system_burst_17 : niosII_system_burst_17
    port map(
      reg_downstream_address => niosII_system_burst_17_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_17_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_17_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_17_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_17_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_17_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_17_downstream_read,
      reg_downstream_write => niosII_system_burst_17_downstream_write,
      reg_downstream_writedata => niosII_system_burst_17_downstream_writedata,
      upstream_readdata => niosII_system_burst_17_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_17_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_17_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_17_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_17_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_17_downstream_waitrequest,
      reset_n => niosII_system_burst_17_downstream_reset_n,
      upstream_address => niosII_system_burst_17_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_17_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_17_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_17_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_17_upstream_address,
      upstream_read => niosII_system_burst_17_upstream_read,
      upstream_write => niosII_system_burst_17_upstream_write,
      upstream_writedata => niosII_system_burst_17_upstream_writedata
    );


  --the_niosII_system_burst_18_upstream, which is an e_instance
  the_niosII_system_burst_18_upstream : niosII_system_burst_18_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_18_upstream => cpu_data_master_granted_niosII_system_burst_18_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_18_upstream => cpu_data_master_qualified_request_niosII_system_burst_18_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_18_upstream => cpu_data_master_requests_niosII_system_burst_18_upstream,
      d1_niosII_system_burst_18_upstream_end_xfer => d1_niosII_system_burst_18_upstream_end_xfer,
      niosII_system_burst_18_upstream_address => niosII_system_burst_18_upstream_address,
      niosII_system_burst_18_upstream_burstcount => niosII_system_burst_18_upstream_burstcount,
      niosII_system_burst_18_upstream_byteaddress => niosII_system_burst_18_upstream_byteaddress,
      niosII_system_burst_18_upstream_byteenable => niosII_system_burst_18_upstream_byteenable,
      niosII_system_burst_18_upstream_debugaccess => niosII_system_burst_18_upstream_debugaccess,
      niosII_system_burst_18_upstream_read => niosII_system_burst_18_upstream_read,
      niosII_system_burst_18_upstream_readdata_from_sa => niosII_system_burst_18_upstream_readdata_from_sa,
      niosII_system_burst_18_upstream_waitrequest_from_sa => niosII_system_burst_18_upstream_waitrequest_from_sa,
      niosII_system_burst_18_upstream_write => niosII_system_burst_18_upstream_write,
      niosII_system_burst_18_upstream_writedata => niosII_system_burst_18_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_18_upstream_readdata => niosII_system_burst_18_upstream_readdata,
      niosII_system_burst_18_upstream_readdatavalid => niosII_system_burst_18_upstream_readdatavalid,
      niosII_system_burst_18_upstream_waitrequest => niosII_system_burst_18_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_18_downstream, which is an e_instance
  the_niosII_system_burst_18_downstream : niosII_system_burst_18_downstream_arbitrator
    port map(
      niosII_system_burst_18_downstream_address_to_slave => niosII_system_burst_18_downstream_address_to_slave,
      niosII_system_burst_18_downstream_latency_counter => niosII_system_burst_18_downstream_latency_counter,
      niosII_system_burst_18_downstream_readdata => niosII_system_burst_18_downstream_readdata,
      niosII_system_burst_18_downstream_readdatavalid => niosII_system_burst_18_downstream_readdatavalid,
      niosII_system_burst_18_downstream_reset_n => niosII_system_burst_18_downstream_reset_n,
      niosII_system_burst_18_downstream_waitrequest => niosII_system_burst_18_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_uart_1_s1_end_xfer => d1_uart_1_s1_end_xfer,
      niosII_system_burst_18_downstream_address => niosII_system_burst_18_downstream_address,
      niosII_system_burst_18_downstream_burstcount => niosII_system_burst_18_downstream_burstcount,
      niosII_system_burst_18_downstream_byteenable => niosII_system_burst_18_downstream_byteenable,
      niosII_system_burst_18_downstream_granted_uart_1_s1 => niosII_system_burst_18_downstream_granted_uart_1_s1,
      niosII_system_burst_18_downstream_qualified_request_uart_1_s1 => niosII_system_burst_18_downstream_qualified_request_uart_1_s1,
      niosII_system_burst_18_downstream_read => niosII_system_burst_18_downstream_read,
      niosII_system_burst_18_downstream_read_data_valid_uart_1_s1 => niosII_system_burst_18_downstream_read_data_valid_uart_1_s1,
      niosII_system_burst_18_downstream_requests_uart_1_s1 => niosII_system_burst_18_downstream_requests_uart_1_s1,
      niosII_system_burst_18_downstream_write => niosII_system_burst_18_downstream_write,
      niosII_system_burst_18_downstream_writedata => niosII_system_burst_18_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      uart_1_s1_readdata_from_sa => uart_1_s1_readdata_from_sa
    );


  --the_niosII_system_burst_18, which is an e_ptf_instance
  the_niosII_system_burst_18 : niosII_system_burst_18
    port map(
      reg_downstream_address => niosII_system_burst_18_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_18_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_18_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_18_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_18_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_18_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_18_downstream_read,
      reg_downstream_write => niosII_system_burst_18_downstream_write,
      reg_downstream_writedata => niosII_system_burst_18_downstream_writedata,
      upstream_readdata => niosII_system_burst_18_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_18_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_18_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_18_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_18_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_18_downstream_waitrequest,
      reset_n => niosII_system_burst_18_downstream_reset_n,
      upstream_address => niosII_system_burst_18_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_18_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_18_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_18_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_18_upstream_address,
      upstream_read => niosII_system_burst_18_upstream_read,
      upstream_write => niosII_system_burst_18_upstream_write,
      upstream_writedata => niosII_system_burst_18_upstream_writedata
    );


  --the_niosII_system_burst_19_upstream, which is an e_instance
  the_niosII_system_burst_19_upstream : niosII_system_burst_19_upstream_arbitrator
    port map(
      cpu_instruction_master_granted_niosII_system_burst_19_upstream => cpu_instruction_master_granted_niosII_system_burst_19_upstream,
      cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream => cpu_instruction_master_qualified_request_niosII_system_burst_19_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream => cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register,
      cpu_instruction_master_requests_niosII_system_burst_19_upstream => cpu_instruction_master_requests_niosII_system_burst_19_upstream,
      d1_niosII_system_burst_19_upstream_end_xfer => d1_niosII_system_burst_19_upstream_end_xfer,
      niosII_system_burst_19_upstream_address => niosII_system_burst_19_upstream_address,
      niosII_system_burst_19_upstream_byteaddress => niosII_system_burst_19_upstream_byteaddress,
      niosII_system_burst_19_upstream_byteenable => niosII_system_burst_19_upstream_byteenable,
      niosII_system_burst_19_upstream_debugaccess => niosII_system_burst_19_upstream_debugaccess,
      niosII_system_burst_19_upstream_read => niosII_system_burst_19_upstream_read,
      niosII_system_burst_19_upstream_readdata_from_sa => niosII_system_burst_19_upstream_readdata_from_sa,
      niosII_system_burst_19_upstream_waitrequest_from_sa => niosII_system_burst_19_upstream_waitrequest_from_sa,
      niosII_system_burst_19_upstream_write => niosII_system_burst_19_upstream_write,
      clk => internal_altpll_inst_c1_out,
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_burstcount => cpu_instruction_master_burstcount,
      cpu_instruction_master_dbs_address => cpu_instruction_master_dbs_address,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register,
      niosII_system_burst_19_upstream_readdata => niosII_system_burst_19_upstream_readdata,
      niosII_system_burst_19_upstream_readdatavalid => niosII_system_burst_19_upstream_readdatavalid,
      niosII_system_burst_19_upstream_waitrequest => niosII_system_burst_19_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_19_downstream, which is an e_instance
  the_niosII_system_burst_19_downstream : niosII_system_burst_19_downstream_arbitrator
    port map(
      niosII_system_burst_19_downstream_address_to_slave => niosII_system_burst_19_downstream_address_to_slave,
      niosII_system_burst_19_downstream_latency_counter => niosII_system_burst_19_downstream_latency_counter,
      niosII_system_burst_19_downstream_readdata => niosII_system_burst_19_downstream_readdata,
      niosII_system_burst_19_downstream_readdatavalid => niosII_system_burst_19_downstream_readdatavalid,
      niosII_system_burst_19_downstream_reset_n => niosII_system_burst_19_downstream_reset_n,
      niosII_system_burst_19_downstream_waitrequest => niosII_system_burst_19_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_tsb_avalon_slave_end_xfer => d1_tsb_avalon_slave_end_xfer,
      incoming_sram_IF_0_tsb_data => incoming_sram_IF_0_tsb_data,
      niosII_system_burst_19_downstream_address => niosII_system_burst_19_downstream_address,
      niosII_system_burst_19_downstream_burstcount => niosII_system_burst_19_downstream_burstcount,
      niosII_system_burst_19_downstream_byteenable => niosII_system_burst_19_downstream_byteenable,
      niosII_system_burst_19_downstream_granted_sram_IF_0_tsb => niosII_system_burst_19_downstream_granted_sram_IF_0_tsb,
      niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb => niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb,
      niosII_system_burst_19_downstream_read => niosII_system_burst_19_downstream_read,
      niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb => niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb,
      niosII_system_burst_19_downstream_requests_sram_IF_0_tsb => niosII_system_burst_19_downstream_requests_sram_IF_0_tsb,
      niosII_system_burst_19_downstream_write => niosII_system_burst_19_downstream_write,
      niosII_system_burst_19_downstream_writedata => niosII_system_burst_19_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_19, which is an e_ptf_instance
  the_niosII_system_burst_19 : niosII_system_burst_19
    port map(
      reg_downstream_address => niosII_system_burst_19_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_19_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_19_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_19_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_19_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_19_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_19_downstream_read,
      reg_downstream_write => niosII_system_burst_19_downstream_write,
      reg_downstream_writedata => niosII_system_burst_19_downstream_writedata,
      upstream_readdata => niosII_system_burst_19_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_19_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_19_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_19_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_19_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_19_downstream_waitrequest,
      reset_n => niosII_system_burst_19_downstream_reset_n,
      upstream_address => niosII_system_burst_19_upstream_byteaddress,
      upstream_byteenable => niosII_system_burst_19_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_19_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_19_upstream_address,
      upstream_read => niosII_system_burst_19_upstream_read,
      upstream_write => niosII_system_burst_19_upstream_write,
      upstream_writedata => niosII_system_burst_19_upstream_writedata
    );


  --the_niosII_system_burst_2_upstream, which is an e_instance
  the_niosII_system_burst_2_upstream : niosII_system_burst_2_upstream_arbitrator
    port map(
      cpu_instruction_master_granted_niosII_system_burst_2_upstream => cpu_instruction_master_granted_niosII_system_burst_2_upstream,
      cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream => cpu_instruction_master_qualified_request_niosII_system_burst_2_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream => cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream,
      cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_2_upstream_shift_register,
      cpu_instruction_master_requests_niosII_system_burst_2_upstream => cpu_instruction_master_requests_niosII_system_burst_2_upstream,
      d1_niosII_system_burst_2_upstream_end_xfer => d1_niosII_system_burst_2_upstream_end_xfer,
      niosII_system_burst_2_upstream_address => niosII_system_burst_2_upstream_address,
      niosII_system_burst_2_upstream_byteaddress => niosII_system_burst_2_upstream_byteaddress,
      niosII_system_burst_2_upstream_byteenable => niosII_system_burst_2_upstream_byteenable,
      niosII_system_burst_2_upstream_debugaccess => niosII_system_burst_2_upstream_debugaccess,
      niosII_system_burst_2_upstream_read => niosII_system_burst_2_upstream_read,
      niosII_system_burst_2_upstream_readdata_from_sa => niosII_system_burst_2_upstream_readdata_from_sa,
      niosII_system_burst_2_upstream_waitrequest_from_sa => niosII_system_burst_2_upstream_waitrequest_from_sa,
      niosII_system_burst_2_upstream_write => niosII_system_burst_2_upstream_write,
      clk => internal_altpll_inst_c1_out,
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_burstcount => cpu_instruction_master_burstcount,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_0_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_10_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_12_upstream_shift_register,
      cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register => cpu_instruction_master_read_data_valid_niosII_system_burst_19_upstream_shift_register,
      niosII_system_burst_2_upstream_readdata => niosII_system_burst_2_upstream_readdata,
      niosII_system_burst_2_upstream_readdatavalid => niosII_system_burst_2_upstream_readdatavalid,
      niosII_system_burst_2_upstream_waitrequest => niosII_system_burst_2_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_2_downstream, which is an e_instance
  the_niosII_system_burst_2_downstream : niosII_system_burst_2_downstream_arbitrator
    port map(
      niosII_system_burst_2_downstream_address_to_slave => niosII_system_burst_2_downstream_address_to_slave,
      niosII_system_burst_2_downstream_latency_counter => niosII_system_burst_2_downstream_latency_counter,
      niosII_system_burst_2_downstream_readdata => niosII_system_burst_2_downstream_readdata,
      niosII_system_burst_2_downstream_readdatavalid => niosII_system_burst_2_downstream_readdatavalid,
      niosII_system_burst_2_downstream_reset_n => niosII_system_burst_2_downstream_reset_n,
      niosII_system_burst_2_downstream_waitrequest => niosII_system_burst_2_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_memory_s1_end_xfer => d1_memory_s1_end_xfer,
      memory_s1_readdata_from_sa => memory_s1_readdata_from_sa,
      niosII_system_burst_2_downstream_address => niosII_system_burst_2_downstream_address,
      niosII_system_burst_2_downstream_burstcount => niosII_system_burst_2_downstream_burstcount,
      niosII_system_burst_2_downstream_byteenable => niosII_system_burst_2_downstream_byteenable,
      niosII_system_burst_2_downstream_granted_memory_s1 => niosII_system_burst_2_downstream_granted_memory_s1,
      niosII_system_burst_2_downstream_qualified_request_memory_s1 => niosII_system_burst_2_downstream_qualified_request_memory_s1,
      niosII_system_burst_2_downstream_read => niosII_system_burst_2_downstream_read,
      niosII_system_burst_2_downstream_read_data_valid_memory_s1 => niosII_system_burst_2_downstream_read_data_valid_memory_s1,
      niosII_system_burst_2_downstream_requests_memory_s1 => niosII_system_burst_2_downstream_requests_memory_s1,
      niosII_system_burst_2_downstream_write => niosII_system_burst_2_downstream_write,
      niosII_system_burst_2_downstream_writedata => niosII_system_burst_2_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_2, which is an e_ptf_instance
  the_niosII_system_burst_2 : niosII_system_burst_2
    port map(
      reg_downstream_address => niosII_system_burst_2_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_2_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_2_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_2_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_2_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_2_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_2_downstream_read,
      reg_downstream_write => niosII_system_burst_2_downstream_write,
      reg_downstream_writedata => niosII_system_burst_2_downstream_writedata,
      upstream_readdata => niosII_system_burst_2_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_2_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_2_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_2_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_2_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_2_downstream_waitrequest,
      reset_n => niosII_system_burst_2_downstream_reset_n,
      upstream_address => niosII_system_burst_2_upstream_byteaddress,
      upstream_byteenable => niosII_system_burst_2_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_2_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_2_upstream_address,
      upstream_read => niosII_system_burst_2_upstream_read,
      upstream_write => niosII_system_burst_2_upstream_write,
      upstream_writedata => niosII_system_burst_2_upstream_writedata
    );


  --the_niosII_system_burst_20_upstream, which is an e_instance
  the_niosII_system_burst_20_upstream : niosII_system_burst_20_upstream_arbitrator
    port map(
      cpu_data_master_byteenable_niosII_system_burst_20_upstream => cpu_data_master_byteenable_niosII_system_burst_20_upstream,
      cpu_data_master_granted_niosII_system_burst_20_upstream => cpu_data_master_granted_niosII_system_burst_20_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_20_upstream => cpu_data_master_qualified_request_niosII_system_burst_20_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_20_upstream => cpu_data_master_requests_niosII_system_burst_20_upstream,
      d1_niosII_system_burst_20_upstream_end_xfer => d1_niosII_system_burst_20_upstream_end_xfer,
      niosII_system_burst_20_upstream_address => niosII_system_burst_20_upstream_address,
      niosII_system_burst_20_upstream_burstcount => niosII_system_burst_20_upstream_burstcount,
      niosII_system_burst_20_upstream_byteaddress => niosII_system_burst_20_upstream_byteaddress,
      niosII_system_burst_20_upstream_byteenable => niosII_system_burst_20_upstream_byteenable,
      niosII_system_burst_20_upstream_debugaccess => niosII_system_burst_20_upstream_debugaccess,
      niosII_system_burst_20_upstream_read => niosII_system_burst_20_upstream_read,
      niosII_system_burst_20_upstream_readdata_from_sa => niosII_system_burst_20_upstream_readdata_from_sa,
      niosII_system_burst_20_upstream_waitrequest_from_sa => niosII_system_burst_20_upstream_waitrequest_from_sa,
      niosII_system_burst_20_upstream_write => niosII_system_burst_20_upstream_write,
      niosII_system_burst_20_upstream_writedata => niosII_system_burst_20_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_dbs_address => cpu_data_master_dbs_address,
      cpu_data_master_dbs_write_16 => cpu_data_master_dbs_write_16,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      niosII_system_burst_20_upstream_readdata => niosII_system_burst_20_upstream_readdata,
      niosII_system_burst_20_upstream_readdatavalid => niosII_system_burst_20_upstream_readdatavalid,
      niosII_system_burst_20_upstream_waitrequest => niosII_system_burst_20_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_20_downstream, which is an e_instance
  the_niosII_system_burst_20_downstream : niosII_system_burst_20_downstream_arbitrator
    port map(
      niosII_system_burst_20_downstream_address_to_slave => niosII_system_burst_20_downstream_address_to_slave,
      niosII_system_burst_20_downstream_latency_counter => niosII_system_burst_20_downstream_latency_counter,
      niosII_system_burst_20_downstream_readdata => niosII_system_burst_20_downstream_readdata,
      niosII_system_burst_20_downstream_readdatavalid => niosII_system_burst_20_downstream_readdatavalid,
      niosII_system_burst_20_downstream_reset_n => niosII_system_burst_20_downstream_reset_n,
      niosII_system_burst_20_downstream_waitrequest => niosII_system_burst_20_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_tsb_avalon_slave_end_xfer => d1_tsb_avalon_slave_end_xfer,
      incoming_sram_IF_0_tsb_data => incoming_sram_IF_0_tsb_data,
      niosII_system_burst_20_downstream_address => niosII_system_burst_20_downstream_address,
      niosII_system_burst_20_downstream_burstcount => niosII_system_burst_20_downstream_burstcount,
      niosII_system_burst_20_downstream_byteenable => niosII_system_burst_20_downstream_byteenable,
      niosII_system_burst_20_downstream_granted_sram_IF_0_tsb => niosII_system_burst_20_downstream_granted_sram_IF_0_tsb,
      niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb => niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb,
      niosII_system_burst_20_downstream_read => niosII_system_burst_20_downstream_read,
      niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb => niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb,
      niosII_system_burst_20_downstream_requests_sram_IF_0_tsb => niosII_system_burst_20_downstream_requests_sram_IF_0_tsb,
      niosII_system_burst_20_downstream_write => niosII_system_burst_20_downstream_write,
      niosII_system_burst_20_downstream_writedata => niosII_system_burst_20_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_20, which is an e_ptf_instance
  the_niosII_system_burst_20 : niosII_system_burst_20
    port map(
      reg_downstream_address => niosII_system_burst_20_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_20_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_20_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_20_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_20_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_20_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_20_downstream_read,
      reg_downstream_write => niosII_system_burst_20_downstream_write,
      reg_downstream_writedata => niosII_system_burst_20_downstream_writedata,
      upstream_readdata => niosII_system_burst_20_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_20_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_20_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_20_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_20_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_20_downstream_waitrequest,
      reset_n => niosII_system_burst_20_downstream_reset_n,
      upstream_address => niosII_system_burst_20_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_20_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_20_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_20_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_20_upstream_address,
      upstream_read => niosII_system_burst_20_upstream_read,
      upstream_write => niosII_system_burst_20_upstream_write,
      upstream_writedata => niosII_system_burst_20_upstream_writedata
    );


  --the_niosII_system_burst_21_upstream, which is an e_instance
  the_niosII_system_burst_21_upstream : niosII_system_burst_21_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_21_upstream => cpu_data_master_granted_niosII_system_burst_21_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_21_upstream => cpu_data_master_qualified_request_niosII_system_burst_21_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_21_upstream => cpu_data_master_requests_niosII_system_burst_21_upstream,
      d1_niosII_system_burst_21_upstream_end_xfer => d1_niosII_system_burst_21_upstream_end_xfer,
      niosII_system_burst_21_upstream_address => niosII_system_burst_21_upstream_address,
      niosII_system_burst_21_upstream_burstcount => niosII_system_burst_21_upstream_burstcount,
      niosII_system_burst_21_upstream_byteaddress => niosII_system_burst_21_upstream_byteaddress,
      niosII_system_burst_21_upstream_byteenable => niosII_system_burst_21_upstream_byteenable,
      niosII_system_burst_21_upstream_debugaccess => niosII_system_burst_21_upstream_debugaccess,
      niosII_system_burst_21_upstream_read => niosII_system_burst_21_upstream_read,
      niosII_system_burst_21_upstream_readdata_from_sa => niosII_system_burst_21_upstream_readdata_from_sa,
      niosII_system_burst_21_upstream_waitrequest_from_sa => niosII_system_burst_21_upstream_waitrequest_from_sa,
      niosII_system_burst_21_upstream_write => niosII_system_burst_21_upstream_write,
      niosII_system_burst_21_upstream_writedata => niosII_system_burst_21_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_21_upstream_readdata => niosII_system_burst_21_upstream_readdata,
      niosII_system_burst_21_upstream_readdatavalid => niosII_system_burst_21_upstream_readdatavalid,
      niosII_system_burst_21_upstream_waitrequest => niosII_system_burst_21_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_21_downstream, which is an e_instance
  the_niosII_system_burst_21_downstream : niosII_system_burst_21_downstream_arbitrator
    port map(
      niosII_system_burst_21_downstream_address_to_slave => niosII_system_burst_21_downstream_address_to_slave,
      niosII_system_burst_21_downstream_latency_counter => niosII_system_burst_21_downstream_latency_counter,
      niosII_system_burst_21_downstream_readdata => niosII_system_burst_21_downstream_readdata,
      niosII_system_burst_21_downstream_readdatavalid => niosII_system_burst_21_downstream_readdatavalid,
      niosII_system_burst_21_downstream_reset_n => niosII_system_burst_21_downstream_reset_n,
      niosII_system_burst_21_downstream_waitrequest => niosII_system_burst_21_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_niosII_system_clock_0_in_end_xfer => d1_niosII_system_clock_0_in_end_xfer,
      niosII_system_burst_21_downstream_address => niosII_system_burst_21_downstream_address,
      niosII_system_burst_21_downstream_burstcount => niosII_system_burst_21_downstream_burstcount,
      niosII_system_burst_21_downstream_byteenable => niosII_system_burst_21_downstream_byteenable,
      niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in => niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in,
      niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in => niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in,
      niosII_system_burst_21_downstream_read => niosII_system_burst_21_downstream_read,
      niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in => niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in,
      niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in => niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in,
      niosII_system_burst_21_downstream_write => niosII_system_burst_21_downstream_write,
      niosII_system_burst_21_downstream_writedata => niosII_system_burst_21_downstream_writedata,
      niosII_system_clock_0_in_readdata_from_sa => niosII_system_clock_0_in_readdata_from_sa,
      niosII_system_clock_0_in_waitrequest_from_sa => niosII_system_clock_0_in_waitrequest_from_sa,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_21, which is an e_ptf_instance
  the_niosII_system_burst_21 : niosII_system_burst_21
    port map(
      reg_downstream_address => niosII_system_burst_21_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_21_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_21_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_21_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_21_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_21_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_21_downstream_read,
      reg_downstream_write => niosII_system_burst_21_downstream_write,
      reg_downstream_writedata => niosII_system_burst_21_downstream_writedata,
      upstream_readdata => niosII_system_burst_21_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_21_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_21_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_21_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_21_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_21_downstream_waitrequest,
      reset_n => niosII_system_burst_21_downstream_reset_n,
      upstream_address => niosII_system_burst_21_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_21_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_21_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_21_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_21_upstream_address,
      upstream_read => niosII_system_burst_21_upstream_read,
      upstream_write => niosII_system_burst_21_upstream_write,
      upstream_writedata => niosII_system_burst_21_upstream_writedata
    );


  --the_niosII_system_burst_3_upstream, which is an e_instance
  the_niosII_system_burst_3_upstream : niosII_system_burst_3_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_3_upstream => cpu_data_master_granted_niosII_system_burst_3_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_3_upstream => cpu_data_master_qualified_request_niosII_system_burst_3_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_3_upstream => cpu_data_master_requests_niosII_system_burst_3_upstream,
      d1_niosII_system_burst_3_upstream_end_xfer => d1_niosII_system_burst_3_upstream_end_xfer,
      niosII_system_burst_3_upstream_address => niosII_system_burst_3_upstream_address,
      niosII_system_burst_3_upstream_burstcount => niosII_system_burst_3_upstream_burstcount,
      niosII_system_burst_3_upstream_byteaddress => niosII_system_burst_3_upstream_byteaddress,
      niosII_system_burst_3_upstream_byteenable => niosII_system_burst_3_upstream_byteenable,
      niosII_system_burst_3_upstream_debugaccess => niosII_system_burst_3_upstream_debugaccess,
      niosII_system_burst_3_upstream_read => niosII_system_burst_3_upstream_read,
      niosII_system_burst_3_upstream_readdata_from_sa => niosII_system_burst_3_upstream_readdata_from_sa,
      niosII_system_burst_3_upstream_waitrequest_from_sa => niosII_system_burst_3_upstream_waitrequest_from_sa,
      niosII_system_burst_3_upstream_write => niosII_system_burst_3_upstream_write,
      niosII_system_burst_3_upstream_writedata => niosII_system_burst_3_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_3_upstream_readdata => niosII_system_burst_3_upstream_readdata,
      niosII_system_burst_3_upstream_readdatavalid => niosII_system_burst_3_upstream_readdatavalid,
      niosII_system_burst_3_upstream_waitrequest => niosII_system_burst_3_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_3_downstream, which is an e_instance
  the_niosII_system_burst_3_downstream : niosII_system_burst_3_downstream_arbitrator
    port map(
      niosII_system_burst_3_downstream_address_to_slave => niosII_system_burst_3_downstream_address_to_slave,
      niosII_system_burst_3_downstream_latency_counter => niosII_system_burst_3_downstream_latency_counter,
      niosII_system_burst_3_downstream_readdata => niosII_system_burst_3_downstream_readdata,
      niosII_system_burst_3_downstream_readdatavalid => niosII_system_burst_3_downstream_readdatavalid,
      niosII_system_burst_3_downstream_reset_n => niosII_system_burst_3_downstream_reset_n,
      niosII_system_burst_3_downstream_waitrequest => niosII_system_burst_3_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_memory_s1_end_xfer => d1_memory_s1_end_xfer,
      memory_s1_readdata_from_sa => memory_s1_readdata_from_sa,
      niosII_system_burst_3_downstream_address => niosII_system_burst_3_downstream_address,
      niosII_system_burst_3_downstream_burstcount => niosII_system_burst_3_downstream_burstcount,
      niosII_system_burst_3_downstream_byteenable => niosII_system_burst_3_downstream_byteenable,
      niosII_system_burst_3_downstream_granted_memory_s1 => niosII_system_burst_3_downstream_granted_memory_s1,
      niosII_system_burst_3_downstream_qualified_request_memory_s1 => niosII_system_burst_3_downstream_qualified_request_memory_s1,
      niosII_system_burst_3_downstream_read => niosII_system_burst_3_downstream_read,
      niosII_system_burst_3_downstream_read_data_valid_memory_s1 => niosII_system_burst_3_downstream_read_data_valid_memory_s1,
      niosII_system_burst_3_downstream_requests_memory_s1 => niosII_system_burst_3_downstream_requests_memory_s1,
      niosII_system_burst_3_downstream_write => niosII_system_burst_3_downstream_write,
      niosII_system_burst_3_downstream_writedata => niosII_system_burst_3_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_3, which is an e_ptf_instance
  the_niosII_system_burst_3 : niosII_system_burst_3
    port map(
      reg_downstream_address => niosII_system_burst_3_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_3_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_3_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_3_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_3_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_3_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_3_downstream_read,
      reg_downstream_write => niosII_system_burst_3_downstream_write,
      reg_downstream_writedata => niosII_system_burst_3_downstream_writedata,
      upstream_readdata => niosII_system_burst_3_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_3_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_3_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_3_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_3_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_3_downstream_waitrequest,
      reset_n => niosII_system_burst_3_downstream_reset_n,
      upstream_address => niosII_system_burst_3_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_3_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_3_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_3_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_3_upstream_address,
      upstream_read => niosII_system_burst_3_upstream_read,
      upstream_write => niosII_system_burst_3_upstream_write,
      upstream_writedata => niosII_system_burst_3_upstream_writedata
    );


  --the_niosII_system_burst_4_upstream, which is an e_instance
  the_niosII_system_burst_4_upstream : niosII_system_burst_4_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_4_upstream => cpu_data_master_granted_niosII_system_burst_4_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_4_upstream => cpu_data_master_qualified_request_niosII_system_burst_4_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_4_upstream => cpu_data_master_requests_niosII_system_burst_4_upstream,
      d1_niosII_system_burst_4_upstream_end_xfer => d1_niosII_system_burst_4_upstream_end_xfer,
      niosII_system_burst_4_upstream_address => niosII_system_burst_4_upstream_address,
      niosII_system_burst_4_upstream_burstcount => niosII_system_burst_4_upstream_burstcount,
      niosII_system_burst_4_upstream_byteaddress => niosII_system_burst_4_upstream_byteaddress,
      niosII_system_burst_4_upstream_byteenable => niosII_system_burst_4_upstream_byteenable,
      niosII_system_burst_4_upstream_debugaccess => niosII_system_burst_4_upstream_debugaccess,
      niosII_system_burst_4_upstream_read => niosII_system_burst_4_upstream_read,
      niosII_system_burst_4_upstream_readdata_from_sa => niosII_system_burst_4_upstream_readdata_from_sa,
      niosII_system_burst_4_upstream_waitrequest_from_sa => niosII_system_burst_4_upstream_waitrequest_from_sa,
      niosII_system_burst_4_upstream_write => niosII_system_burst_4_upstream_write,
      niosII_system_burst_4_upstream_writedata => niosII_system_burst_4_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_4_upstream_readdata => niosII_system_burst_4_upstream_readdata,
      niosII_system_burst_4_upstream_readdatavalid => niosII_system_burst_4_upstream_readdatavalid,
      niosII_system_burst_4_upstream_waitrequest => niosII_system_burst_4_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_4_downstream, which is an e_instance
  the_niosII_system_burst_4_downstream : niosII_system_burst_4_downstream_arbitrator
    port map(
      niosII_system_burst_4_downstream_address_to_slave => niosII_system_burst_4_downstream_address_to_slave,
      niosII_system_burst_4_downstream_latency_counter => niosII_system_burst_4_downstream_latency_counter,
      niosII_system_burst_4_downstream_readdata => niosII_system_burst_4_downstream_readdata,
      niosII_system_burst_4_downstream_readdatavalid => niosII_system_burst_4_downstream_readdatavalid,
      niosII_system_burst_4_downstream_reset_n => niosII_system_burst_4_downstream_reset_n,
      niosII_system_burst_4_downstream_waitrequest => niosII_system_burst_4_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      niosII_system_burst_4_downstream_address => niosII_system_burst_4_downstream_address,
      niosII_system_burst_4_downstream_burstcount => niosII_system_burst_4_downstream_burstcount,
      niosII_system_burst_4_downstream_byteenable => niosII_system_burst_4_downstream_byteenable,
      niosII_system_burst_4_downstream_granted_sysid_control_slave => niosII_system_burst_4_downstream_granted_sysid_control_slave,
      niosII_system_burst_4_downstream_qualified_request_sysid_control_slave => niosII_system_burst_4_downstream_qualified_request_sysid_control_slave,
      niosII_system_burst_4_downstream_read => niosII_system_burst_4_downstream_read,
      niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave => niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave,
      niosII_system_burst_4_downstream_requests_sysid_control_slave => niosII_system_burst_4_downstream_requests_sysid_control_slave,
      niosII_system_burst_4_downstream_write => niosII_system_burst_4_downstream_write,
      niosII_system_burst_4_downstream_writedata => niosII_system_burst_4_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa
    );


  --the_niosII_system_burst_4, which is an e_ptf_instance
  the_niosII_system_burst_4 : niosII_system_burst_4
    port map(
      reg_downstream_address => niosII_system_burst_4_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_4_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_4_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_4_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_4_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_4_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_4_downstream_read,
      reg_downstream_write => niosII_system_burst_4_downstream_write,
      reg_downstream_writedata => niosII_system_burst_4_downstream_writedata,
      upstream_readdata => niosII_system_burst_4_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_4_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_4_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_4_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_4_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_4_downstream_waitrequest,
      reset_n => niosII_system_burst_4_downstream_reset_n,
      upstream_address => niosII_system_burst_4_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_4_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_4_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_4_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_4_upstream_address,
      upstream_read => niosII_system_burst_4_upstream_read,
      upstream_write => niosII_system_burst_4_upstream_write,
      upstream_writedata => niosII_system_burst_4_upstream_writedata
    );


  --the_niosII_system_burst_5_upstream, which is an e_instance
  the_niosII_system_burst_5_upstream : niosII_system_burst_5_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_5_upstream => cpu_data_master_granted_niosII_system_burst_5_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_5_upstream => cpu_data_master_qualified_request_niosII_system_burst_5_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_5_upstream => cpu_data_master_requests_niosII_system_burst_5_upstream,
      d1_niosII_system_burst_5_upstream_end_xfer => d1_niosII_system_burst_5_upstream_end_xfer,
      niosII_system_burst_5_upstream_address => niosII_system_burst_5_upstream_address,
      niosII_system_burst_5_upstream_burstcount => niosII_system_burst_5_upstream_burstcount,
      niosII_system_burst_5_upstream_byteaddress => niosII_system_burst_5_upstream_byteaddress,
      niosII_system_burst_5_upstream_byteenable => niosII_system_burst_5_upstream_byteenable,
      niosII_system_burst_5_upstream_debugaccess => niosII_system_burst_5_upstream_debugaccess,
      niosII_system_burst_5_upstream_read => niosII_system_burst_5_upstream_read,
      niosII_system_burst_5_upstream_readdata_from_sa => niosII_system_burst_5_upstream_readdata_from_sa,
      niosII_system_burst_5_upstream_waitrequest_from_sa => niosII_system_burst_5_upstream_waitrequest_from_sa,
      niosII_system_burst_5_upstream_write => niosII_system_burst_5_upstream_write,
      niosII_system_burst_5_upstream_writedata => niosII_system_burst_5_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_5_upstream_readdata => niosII_system_burst_5_upstream_readdata,
      niosII_system_burst_5_upstream_readdatavalid => niosII_system_burst_5_upstream_readdatavalid,
      niosII_system_burst_5_upstream_waitrequest => niosII_system_burst_5_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_5_downstream, which is an e_instance
  the_niosII_system_burst_5_downstream : niosII_system_burst_5_downstream_arbitrator
    port map(
      niosII_system_burst_5_downstream_address_to_slave => niosII_system_burst_5_downstream_address_to_slave,
      niosII_system_burst_5_downstream_latency_counter => niosII_system_burst_5_downstream_latency_counter,
      niosII_system_burst_5_downstream_readdata => niosII_system_burst_5_downstream_readdata,
      niosII_system_burst_5_downstream_readdatavalid => niosII_system_burst_5_downstream_readdatavalid,
      niosII_system_burst_5_downstream_reset_n => niosII_system_burst_5_downstream_reset_n,
      niosII_system_burst_5_downstream_waitrequest => niosII_system_burst_5_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_sys_clk_timer_s1_end_xfer => d1_sys_clk_timer_s1_end_xfer,
      niosII_system_burst_5_downstream_address => niosII_system_burst_5_downstream_address,
      niosII_system_burst_5_downstream_burstcount => niosII_system_burst_5_downstream_burstcount,
      niosII_system_burst_5_downstream_byteenable => niosII_system_burst_5_downstream_byteenable,
      niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 => niosII_system_burst_5_downstream_granted_sys_clk_timer_s1,
      niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 => niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1,
      niosII_system_burst_5_downstream_read => niosII_system_burst_5_downstream_read,
      niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1 => niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1,
      niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 => niosII_system_burst_5_downstream_requests_sys_clk_timer_s1,
      niosII_system_burst_5_downstream_write => niosII_system_burst_5_downstream_write,
      niosII_system_burst_5_downstream_writedata => niosII_system_burst_5_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      sys_clk_timer_s1_readdata_from_sa => sys_clk_timer_s1_readdata_from_sa
    );


  --the_niosII_system_burst_5, which is an e_ptf_instance
  the_niosII_system_burst_5 : niosII_system_burst_5
    port map(
      reg_downstream_address => niosII_system_burst_5_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_5_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_5_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_5_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_5_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_5_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_5_downstream_read,
      reg_downstream_write => niosII_system_burst_5_downstream_write,
      reg_downstream_writedata => niosII_system_burst_5_downstream_writedata,
      upstream_readdata => niosII_system_burst_5_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_5_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_5_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_5_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_5_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_5_downstream_waitrequest,
      reset_n => niosII_system_burst_5_downstream_reset_n,
      upstream_address => niosII_system_burst_5_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_5_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_5_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_5_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_5_upstream_address,
      upstream_read => niosII_system_burst_5_upstream_read,
      upstream_write => niosII_system_burst_5_upstream_write,
      upstream_writedata => niosII_system_burst_5_upstream_writedata
    );


  --the_niosII_system_burst_6_upstream, which is an e_instance
  the_niosII_system_burst_6_upstream : niosII_system_burst_6_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_6_upstream => cpu_data_master_granted_niosII_system_burst_6_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_6_upstream => cpu_data_master_qualified_request_niosII_system_burst_6_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_6_upstream => cpu_data_master_requests_niosII_system_burst_6_upstream,
      d1_niosII_system_burst_6_upstream_end_xfer => d1_niosII_system_burst_6_upstream_end_xfer,
      niosII_system_burst_6_upstream_address => niosII_system_burst_6_upstream_address,
      niosII_system_burst_6_upstream_burstcount => niosII_system_burst_6_upstream_burstcount,
      niosII_system_burst_6_upstream_byteaddress => niosII_system_burst_6_upstream_byteaddress,
      niosII_system_burst_6_upstream_byteenable => niosII_system_burst_6_upstream_byteenable,
      niosII_system_burst_6_upstream_debugaccess => niosII_system_burst_6_upstream_debugaccess,
      niosII_system_burst_6_upstream_read => niosII_system_burst_6_upstream_read,
      niosII_system_burst_6_upstream_readdata_from_sa => niosII_system_burst_6_upstream_readdata_from_sa,
      niosII_system_burst_6_upstream_waitrequest_from_sa => niosII_system_burst_6_upstream_waitrequest_from_sa,
      niosII_system_burst_6_upstream_write => niosII_system_burst_6_upstream_write,
      niosII_system_burst_6_upstream_writedata => niosII_system_burst_6_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_6_upstream_readdata => niosII_system_burst_6_upstream_readdata,
      niosII_system_burst_6_upstream_readdatavalid => niosII_system_burst_6_upstream_readdatavalid,
      niosII_system_burst_6_upstream_waitrequest => niosII_system_burst_6_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_6_downstream, which is an e_instance
  the_niosII_system_burst_6_downstream : niosII_system_burst_6_downstream_arbitrator
    port map(
      niosII_system_burst_6_downstream_address_to_slave => niosII_system_burst_6_downstream_address_to_slave,
      niosII_system_burst_6_downstream_latency_counter => niosII_system_burst_6_downstream_latency_counter,
      niosII_system_burst_6_downstream_readdata => niosII_system_burst_6_downstream_readdata,
      niosII_system_burst_6_downstream_readdatavalid => niosII_system_burst_6_downstream_readdatavalid,
      niosII_system_burst_6_downstream_reset_n => niosII_system_burst_6_downstream_reset_n,
      niosII_system_burst_6_downstream_waitrequest => niosII_system_burst_6_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      niosII_system_burst_6_downstream_address => niosII_system_burst_6_downstream_address,
      niosII_system_burst_6_downstream_burstcount => niosII_system_burst_6_downstream_burstcount,
      niosII_system_burst_6_downstream_byteenable => niosII_system_burst_6_downstream_byteenable,
      niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave => niosII_system_burst_6_downstream_granted_jtag_uart_avalon_jtag_slave,
      niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave => niosII_system_burst_6_downstream_qualified_request_jtag_uart_avalon_jtag_slave,
      niosII_system_burst_6_downstream_read => niosII_system_burst_6_downstream_read,
      niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave => niosII_system_burst_6_downstream_read_data_valid_jtag_uart_avalon_jtag_slave,
      niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave => niosII_system_burst_6_downstream_requests_jtag_uart_avalon_jtag_slave,
      niosII_system_burst_6_downstream_write => niosII_system_burst_6_downstream_write,
      niosII_system_burst_6_downstream_writedata => niosII_system_burst_6_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_6, which is an e_ptf_instance
  the_niosII_system_burst_6 : niosII_system_burst_6
    port map(
      reg_downstream_address => niosII_system_burst_6_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_6_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_6_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_6_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_6_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_6_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_6_downstream_read,
      reg_downstream_write => niosII_system_burst_6_downstream_write,
      reg_downstream_writedata => niosII_system_burst_6_downstream_writedata,
      upstream_readdata => niosII_system_burst_6_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_6_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_6_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_6_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_6_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_6_downstream_waitrequest,
      reset_n => niosII_system_burst_6_downstream_reset_n,
      upstream_address => niosII_system_burst_6_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_6_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_6_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_6_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_6_upstream_address,
      upstream_read => niosII_system_burst_6_upstream_read,
      upstream_write => niosII_system_burst_6_upstream_write,
      upstream_writedata => niosII_system_burst_6_upstream_writedata
    );


  --the_niosII_system_burst_7_upstream, which is an e_instance
  the_niosII_system_burst_7_upstream : niosII_system_burst_7_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_7_upstream => cpu_data_master_granted_niosII_system_burst_7_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_7_upstream => cpu_data_master_qualified_request_niosII_system_burst_7_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_7_upstream => cpu_data_master_requests_niosII_system_burst_7_upstream,
      d1_niosII_system_burst_7_upstream_end_xfer => d1_niosII_system_burst_7_upstream_end_xfer,
      niosII_system_burst_7_upstream_address => niosII_system_burst_7_upstream_address,
      niosII_system_burst_7_upstream_burstcount => niosII_system_burst_7_upstream_burstcount,
      niosII_system_burst_7_upstream_byteaddress => niosII_system_burst_7_upstream_byteaddress,
      niosII_system_burst_7_upstream_byteenable => niosII_system_burst_7_upstream_byteenable,
      niosII_system_burst_7_upstream_debugaccess => niosII_system_burst_7_upstream_debugaccess,
      niosII_system_burst_7_upstream_read => niosII_system_burst_7_upstream_read,
      niosII_system_burst_7_upstream_readdata_from_sa => niosII_system_burst_7_upstream_readdata_from_sa,
      niosII_system_burst_7_upstream_waitrequest_from_sa => niosII_system_burst_7_upstream_waitrequest_from_sa,
      niosII_system_burst_7_upstream_write => niosII_system_burst_7_upstream_write,
      niosII_system_burst_7_upstream_writedata => niosII_system_burst_7_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_7_upstream_readdata => niosII_system_burst_7_upstream_readdata,
      niosII_system_burst_7_upstream_readdatavalid => niosII_system_burst_7_upstream_readdatavalid,
      niosII_system_burst_7_upstream_waitrequest => niosII_system_burst_7_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_7_downstream, which is an e_instance
  the_niosII_system_burst_7_downstream : niosII_system_burst_7_downstream_arbitrator
    port map(
      niosII_system_burst_7_downstream_address_to_slave => niosII_system_burst_7_downstream_address_to_slave,
      niosII_system_burst_7_downstream_latency_counter => niosII_system_burst_7_downstream_latency_counter,
      niosII_system_burst_7_downstream_readdata => niosII_system_burst_7_downstream_readdata,
      niosII_system_burst_7_downstream_readdatavalid => niosII_system_burst_7_downstream_readdatavalid,
      niosII_system_burst_7_downstream_reset_n => niosII_system_burst_7_downstream_reset_n,
      niosII_system_burst_7_downstream_waitrequest => niosII_system_burst_7_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_lcd_display_control_slave_end_xfer => d1_lcd_display_control_slave_end_xfer,
      lcd_display_control_slave_readdata_from_sa => lcd_display_control_slave_readdata_from_sa,
      lcd_display_control_slave_wait_counter_eq_0 => lcd_display_control_slave_wait_counter_eq_0,
      niosII_system_burst_7_downstream_address => niosII_system_burst_7_downstream_address,
      niosII_system_burst_7_downstream_burstcount => niosII_system_burst_7_downstream_burstcount,
      niosII_system_burst_7_downstream_byteenable => niosII_system_burst_7_downstream_byteenable,
      niosII_system_burst_7_downstream_granted_lcd_display_control_slave => niosII_system_burst_7_downstream_granted_lcd_display_control_slave,
      niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave => niosII_system_burst_7_downstream_qualified_request_lcd_display_control_slave,
      niosII_system_burst_7_downstream_read => niosII_system_burst_7_downstream_read,
      niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave => niosII_system_burst_7_downstream_read_data_valid_lcd_display_control_slave,
      niosII_system_burst_7_downstream_requests_lcd_display_control_slave => niosII_system_burst_7_downstream_requests_lcd_display_control_slave,
      niosII_system_burst_7_downstream_write => niosII_system_burst_7_downstream_write,
      niosII_system_burst_7_downstream_writedata => niosII_system_burst_7_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_7, which is an e_ptf_instance
  the_niosII_system_burst_7 : niosII_system_burst_7
    port map(
      reg_downstream_address => niosII_system_burst_7_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_7_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_7_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_7_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_7_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_7_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_7_downstream_read,
      reg_downstream_write => niosII_system_burst_7_downstream_write,
      reg_downstream_writedata => niosII_system_burst_7_downstream_writedata,
      upstream_readdata => niosII_system_burst_7_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_7_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_7_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_7_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_7_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_7_downstream_waitrequest,
      reset_n => niosII_system_burst_7_downstream_reset_n,
      upstream_address => niosII_system_burst_7_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_7_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_7_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_7_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_7_upstream_address,
      upstream_read => niosII_system_burst_7_upstream_read,
      upstream_write => niosII_system_burst_7_upstream_write,
      upstream_writedata => niosII_system_burst_7_upstream_writedata
    );


  --the_niosII_system_burst_8_upstream, which is an e_instance
  the_niosII_system_burst_8_upstream : niosII_system_burst_8_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_8_upstream => cpu_data_master_granted_niosII_system_burst_8_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_8_upstream => cpu_data_master_qualified_request_niosII_system_burst_8_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_8_upstream => cpu_data_master_requests_niosII_system_burst_8_upstream,
      d1_niosII_system_burst_8_upstream_end_xfer => d1_niosII_system_burst_8_upstream_end_xfer,
      niosII_system_burst_8_upstream_address => niosII_system_burst_8_upstream_address,
      niosII_system_burst_8_upstream_burstcount => niosII_system_burst_8_upstream_burstcount,
      niosII_system_burst_8_upstream_byteaddress => niosII_system_burst_8_upstream_byteaddress,
      niosII_system_burst_8_upstream_byteenable => niosII_system_burst_8_upstream_byteenable,
      niosII_system_burst_8_upstream_debugaccess => niosII_system_burst_8_upstream_debugaccess,
      niosII_system_burst_8_upstream_read => niosII_system_burst_8_upstream_read,
      niosII_system_burst_8_upstream_readdata_from_sa => niosII_system_burst_8_upstream_readdata_from_sa,
      niosII_system_burst_8_upstream_waitrequest_from_sa => niosII_system_burst_8_upstream_waitrequest_from_sa,
      niosII_system_burst_8_upstream_write => niosII_system_burst_8_upstream_write,
      niosII_system_burst_8_upstream_writedata => niosII_system_burst_8_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_8_upstream_readdata => niosII_system_burst_8_upstream_readdata,
      niosII_system_burst_8_upstream_readdatavalid => niosII_system_burst_8_upstream_readdatavalid,
      niosII_system_burst_8_upstream_waitrequest => niosII_system_burst_8_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_8_downstream, which is an e_instance
  the_niosII_system_burst_8_downstream : niosII_system_burst_8_downstream_arbitrator
    port map(
      niosII_system_burst_8_downstream_address_to_slave => niosII_system_burst_8_downstream_address_to_slave,
      niosII_system_burst_8_downstream_latency_counter => niosII_system_burst_8_downstream_latency_counter,
      niosII_system_burst_8_downstream_readdata => niosII_system_burst_8_downstream_readdata,
      niosII_system_burst_8_downstream_readdatavalid => niosII_system_burst_8_downstream_readdatavalid,
      niosII_system_burst_8_downstream_reset_n => niosII_system_burst_8_downstream_reset_n,
      niosII_system_burst_8_downstream_waitrequest => niosII_system_burst_8_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_led_pio_s1_end_xfer => d1_led_pio_s1_end_xfer,
      led_pio_s1_readdata_from_sa => led_pio_s1_readdata_from_sa,
      niosII_system_burst_8_downstream_address => niosII_system_burst_8_downstream_address,
      niosII_system_burst_8_downstream_burstcount => niosII_system_burst_8_downstream_burstcount,
      niosII_system_burst_8_downstream_byteenable => niosII_system_burst_8_downstream_byteenable,
      niosII_system_burst_8_downstream_granted_led_pio_s1 => niosII_system_burst_8_downstream_granted_led_pio_s1,
      niosII_system_burst_8_downstream_qualified_request_led_pio_s1 => niosII_system_burst_8_downstream_qualified_request_led_pio_s1,
      niosII_system_burst_8_downstream_read => niosII_system_burst_8_downstream_read,
      niosII_system_burst_8_downstream_read_data_valid_led_pio_s1 => niosII_system_burst_8_downstream_read_data_valid_led_pio_s1,
      niosII_system_burst_8_downstream_requests_led_pio_s1 => niosII_system_burst_8_downstream_requests_led_pio_s1,
      niosII_system_burst_8_downstream_write => niosII_system_burst_8_downstream_write,
      niosII_system_burst_8_downstream_writedata => niosII_system_burst_8_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_8, which is an e_ptf_instance
  the_niosII_system_burst_8 : niosII_system_burst_8
    port map(
      reg_downstream_address => niosII_system_burst_8_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_8_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_8_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_8_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_8_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_8_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_8_downstream_read,
      reg_downstream_write => niosII_system_burst_8_downstream_write,
      reg_downstream_writedata => niosII_system_burst_8_downstream_writedata,
      upstream_readdata => niosII_system_burst_8_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_8_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_8_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_8_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_8_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_8_downstream_waitrequest,
      reset_n => niosII_system_burst_8_downstream_reset_n,
      upstream_address => niosII_system_burst_8_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_8_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_8_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_8_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_8_upstream_address,
      upstream_read => niosII_system_burst_8_upstream_read,
      upstream_write => niosII_system_burst_8_upstream_write,
      upstream_writedata => niosII_system_burst_8_upstream_writedata
    );


  --the_niosII_system_burst_9_upstream, which is an e_instance
  the_niosII_system_burst_9_upstream : niosII_system_burst_9_upstream_arbitrator
    port map(
      cpu_data_master_granted_niosII_system_burst_9_upstream => cpu_data_master_granted_niosII_system_burst_9_upstream,
      cpu_data_master_qualified_request_niosII_system_burst_9_upstream => cpu_data_master_qualified_request_niosII_system_burst_9_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream,
      cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_9_upstream_shift_register,
      cpu_data_master_requests_niosII_system_burst_9_upstream => cpu_data_master_requests_niosII_system_burst_9_upstream,
      d1_niosII_system_burst_9_upstream_end_xfer => d1_niosII_system_burst_9_upstream_end_xfer,
      niosII_system_burst_9_upstream_address => niosII_system_burst_9_upstream_address,
      niosII_system_burst_9_upstream_burstcount => niosII_system_burst_9_upstream_burstcount,
      niosII_system_burst_9_upstream_byteaddress => niosII_system_burst_9_upstream_byteaddress,
      niosII_system_burst_9_upstream_byteenable => niosII_system_burst_9_upstream_byteenable,
      niosII_system_burst_9_upstream_debugaccess => niosII_system_burst_9_upstream_debugaccess,
      niosII_system_burst_9_upstream_read => niosII_system_burst_9_upstream_read,
      niosII_system_burst_9_upstream_readdata_from_sa => niosII_system_burst_9_upstream_readdata_from_sa,
      niosII_system_burst_9_upstream_waitrequest_from_sa => niosII_system_burst_9_upstream_waitrequest_from_sa,
      niosII_system_burst_9_upstream_write => niosII_system_burst_9_upstream_write,
      niosII_system_burst_9_upstream_writedata => niosII_system_burst_9_upstream_writedata,
      clk => internal_altpll_inst_c1_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_burstcount => cpu_data_master_burstcount,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_11_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_13_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_14_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_15_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_16_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_17_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_18_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_1_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_20_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_21_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_3_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_4_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_5_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_6_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_7_upstream_shift_register,
      cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register => cpu_data_master_read_data_valid_niosII_system_burst_8_upstream_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      niosII_system_burst_9_upstream_readdata => niosII_system_burst_9_upstream_readdata,
      niosII_system_burst_9_upstream_readdatavalid => niosII_system_burst_9_upstream_readdatavalid,
      niosII_system_burst_9_upstream_waitrequest => niosII_system_burst_9_upstream_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_burst_9_downstream, which is an e_instance
  the_niosII_system_burst_9_downstream : niosII_system_burst_9_downstream_arbitrator
    port map(
      niosII_system_burst_9_downstream_address_to_slave => niosII_system_burst_9_downstream_address_to_slave,
      niosII_system_burst_9_downstream_latency_counter => niosII_system_burst_9_downstream_latency_counter,
      niosII_system_burst_9_downstream_readdata => niosII_system_burst_9_downstream_readdata,
      niosII_system_burst_9_downstream_readdatavalid => niosII_system_burst_9_downstream_readdatavalid,
      niosII_system_burst_9_downstream_reset_n => niosII_system_burst_9_downstream_reset_n,
      niosII_system_burst_9_downstream_waitrequest => niosII_system_burst_9_downstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      d1_switch_s1_end_xfer => d1_switch_s1_end_xfer,
      niosII_system_burst_9_downstream_address => niosII_system_burst_9_downstream_address,
      niosII_system_burst_9_downstream_burstcount => niosII_system_burst_9_downstream_burstcount,
      niosII_system_burst_9_downstream_byteenable => niosII_system_burst_9_downstream_byteenable,
      niosII_system_burst_9_downstream_granted_switch_s1 => niosII_system_burst_9_downstream_granted_switch_s1,
      niosII_system_burst_9_downstream_qualified_request_switch_s1 => niosII_system_burst_9_downstream_qualified_request_switch_s1,
      niosII_system_burst_9_downstream_read => niosII_system_burst_9_downstream_read,
      niosII_system_burst_9_downstream_read_data_valid_switch_s1 => niosII_system_burst_9_downstream_read_data_valid_switch_s1,
      niosII_system_burst_9_downstream_requests_switch_s1 => niosII_system_burst_9_downstream_requests_switch_s1,
      niosII_system_burst_9_downstream_write => niosII_system_burst_9_downstream_write,
      niosII_system_burst_9_downstream_writedata => niosII_system_burst_9_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      switch_s1_readdata_from_sa => switch_s1_readdata_from_sa
    );


  --the_niosII_system_burst_9, which is an e_ptf_instance
  the_niosII_system_burst_9 : niosII_system_burst_9
    port map(
      reg_downstream_address => niosII_system_burst_9_downstream_address,
      reg_downstream_arbitrationshare => niosII_system_burst_9_downstream_arbitrationshare,
      reg_downstream_burstcount => niosII_system_burst_9_downstream_burstcount,
      reg_downstream_byteenable => niosII_system_burst_9_downstream_byteenable,
      reg_downstream_debugaccess => niosII_system_burst_9_downstream_debugaccess,
      reg_downstream_nativeaddress => niosII_system_burst_9_downstream_nativeaddress,
      reg_downstream_read => niosII_system_burst_9_downstream_read,
      reg_downstream_write => niosII_system_burst_9_downstream_write,
      reg_downstream_writedata => niosII_system_burst_9_downstream_writedata,
      upstream_readdata => niosII_system_burst_9_upstream_readdata,
      upstream_readdatavalid => niosII_system_burst_9_upstream_readdatavalid,
      upstream_waitrequest => niosII_system_burst_9_upstream_waitrequest,
      clk => internal_altpll_inst_c1_out,
      downstream_readdata => niosII_system_burst_9_downstream_readdata,
      downstream_readdatavalid => niosII_system_burst_9_downstream_readdatavalid,
      downstream_waitrequest => niosII_system_burst_9_downstream_waitrequest,
      reset_n => niosII_system_burst_9_downstream_reset_n,
      upstream_address => niosII_system_burst_9_upstream_byteaddress,
      upstream_burstcount => niosII_system_burst_9_upstream_burstcount,
      upstream_byteenable => niosII_system_burst_9_upstream_byteenable,
      upstream_debugaccess => niosII_system_burst_9_upstream_debugaccess,
      upstream_nativeaddress => niosII_system_burst_9_upstream_address,
      upstream_read => niosII_system_burst_9_upstream_read,
      upstream_write => niosII_system_burst_9_upstream_write,
      upstream_writedata => niosII_system_burst_9_upstream_writedata
    );


  --the_niosII_system_clock_0_in, which is an e_instance
  the_niosII_system_clock_0_in : niosII_system_clock_0_in_arbitrator
    port map(
      d1_niosII_system_clock_0_in_end_xfer => d1_niosII_system_clock_0_in_end_xfer,
      niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in => niosII_system_burst_21_downstream_granted_niosII_system_clock_0_in,
      niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in => niosII_system_burst_21_downstream_qualified_request_niosII_system_clock_0_in,
      niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in => niosII_system_burst_21_downstream_read_data_valid_niosII_system_clock_0_in,
      niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in => niosII_system_burst_21_downstream_requests_niosII_system_clock_0_in,
      niosII_system_clock_0_in_address => niosII_system_clock_0_in_address,
      niosII_system_clock_0_in_byteenable => niosII_system_clock_0_in_byteenable,
      niosII_system_clock_0_in_endofpacket_from_sa => niosII_system_clock_0_in_endofpacket_from_sa,
      niosII_system_clock_0_in_nativeaddress => niosII_system_clock_0_in_nativeaddress,
      niosII_system_clock_0_in_read => niosII_system_clock_0_in_read,
      niosII_system_clock_0_in_readdata_from_sa => niosII_system_clock_0_in_readdata_from_sa,
      niosII_system_clock_0_in_reset_n => niosII_system_clock_0_in_reset_n,
      niosII_system_clock_0_in_waitrequest_from_sa => niosII_system_clock_0_in_waitrequest_from_sa,
      niosII_system_clock_0_in_write => niosII_system_clock_0_in_write,
      niosII_system_clock_0_in_writedata => niosII_system_clock_0_in_writedata,
      clk => internal_altpll_inst_c1_out,
      niosII_system_burst_21_downstream_address_to_slave => niosII_system_burst_21_downstream_address_to_slave,
      niosII_system_burst_21_downstream_arbitrationshare => niosII_system_burst_21_downstream_arbitrationshare,
      niosII_system_burst_21_downstream_burstcount => niosII_system_burst_21_downstream_burstcount,
      niosII_system_burst_21_downstream_byteenable => niosII_system_burst_21_downstream_byteenable,
      niosII_system_burst_21_downstream_latency_counter => niosII_system_burst_21_downstream_latency_counter,
      niosII_system_burst_21_downstream_nativeaddress => niosII_system_burst_21_downstream_nativeaddress,
      niosII_system_burst_21_downstream_read => niosII_system_burst_21_downstream_read,
      niosII_system_burst_21_downstream_write => niosII_system_burst_21_downstream_write,
      niosII_system_burst_21_downstream_writedata => niosII_system_burst_21_downstream_writedata,
      niosII_system_clock_0_in_endofpacket => niosII_system_clock_0_in_endofpacket,
      niosII_system_clock_0_in_readdata => niosII_system_clock_0_in_readdata,
      niosII_system_clock_0_in_waitrequest => niosII_system_clock_0_in_waitrequest,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_niosII_system_clock_0_out, which is an e_instance
  the_niosII_system_clock_0_out : niosII_system_clock_0_out_arbitrator
    port map(
      niosII_system_clock_0_out_address_to_slave => niosII_system_clock_0_out_address_to_slave,
      niosII_system_clock_0_out_readdata => niosII_system_clock_0_out_readdata,
      niosII_system_clock_0_out_reset_n => niosII_system_clock_0_out_reset_n,
      niosII_system_clock_0_out_waitrequest => niosII_system_clock_0_out_waitrequest,
      altpll_inst_pll_slave_readdata_from_sa => altpll_inst_pll_slave_readdata_from_sa,
      clk => clk_0,
      d1_altpll_inst_pll_slave_end_xfer => d1_altpll_inst_pll_slave_end_xfer,
      niosII_system_clock_0_out_address => niosII_system_clock_0_out_address,
      niosII_system_clock_0_out_byteenable => niosII_system_clock_0_out_byteenable,
      niosII_system_clock_0_out_granted_altpll_inst_pll_slave => niosII_system_clock_0_out_granted_altpll_inst_pll_slave,
      niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave => niosII_system_clock_0_out_qualified_request_altpll_inst_pll_slave,
      niosII_system_clock_0_out_read => niosII_system_clock_0_out_read,
      niosII_system_clock_0_out_read_data_valid_altpll_inst_pll_slave => niosII_system_clock_0_out_read_data_valid_altpll_inst_pll_slave,
      niosII_system_clock_0_out_requests_altpll_inst_pll_slave => niosII_system_clock_0_out_requests_altpll_inst_pll_slave,
      niosII_system_clock_0_out_write => niosII_system_clock_0_out_write,
      niosII_system_clock_0_out_writedata => niosII_system_clock_0_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_niosII_system_clock_0, which is an e_ptf_instance
  the_niosII_system_clock_0 : niosII_system_clock_0
    port map(
      master_address => niosII_system_clock_0_out_address,
      master_byteenable => niosII_system_clock_0_out_byteenable,
      master_nativeaddress => niosII_system_clock_0_out_nativeaddress,
      master_read => niosII_system_clock_0_out_read,
      master_write => niosII_system_clock_0_out_write,
      master_writedata => niosII_system_clock_0_out_writedata,
      slave_endofpacket => niosII_system_clock_0_in_endofpacket,
      slave_readdata => niosII_system_clock_0_in_readdata,
      slave_waitrequest => niosII_system_clock_0_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => niosII_system_clock_0_out_endofpacket,
      master_readdata => niosII_system_clock_0_out_readdata,
      master_reset_n => niosII_system_clock_0_out_reset_n,
      master_waitrequest => niosII_system_clock_0_out_waitrequest,
      slave_address => niosII_system_clock_0_in_address,
      slave_byteenable => niosII_system_clock_0_in_byteenable,
      slave_clk => internal_altpll_inst_c1_out,
      slave_nativeaddress => niosII_system_clock_0_in_nativeaddress,
      slave_read => niosII_system_clock_0_in_read,
      slave_reset_n => niosII_system_clock_0_in_reset_n,
      slave_write => niosII_system_clock_0_in_write,
      slave_writedata => niosII_system_clock_0_in_writedata
    );


  --the_sdram_s1, which is an e_instance
  the_sdram_s1 : sdram_s1_arbitrator
    port map(
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      niosII_system_burst_10_downstream_granted_sdram_s1 => niosII_system_burst_10_downstream_granted_sdram_s1,
      niosII_system_burst_10_downstream_qualified_request_sdram_s1 => niosII_system_burst_10_downstream_qualified_request_sdram_s1,
      niosII_system_burst_10_downstream_read_data_valid_sdram_s1 => niosII_system_burst_10_downstream_read_data_valid_sdram_s1,
      niosII_system_burst_10_downstream_read_data_valid_sdram_s1_shift_register => niosII_system_burst_10_downstream_read_data_valid_sdram_s1_shift_register,
      niosII_system_burst_10_downstream_requests_sdram_s1 => niosII_system_burst_10_downstream_requests_sdram_s1,
      niosII_system_burst_11_downstream_granted_sdram_s1 => niosII_system_burst_11_downstream_granted_sdram_s1,
      niosII_system_burst_11_downstream_qualified_request_sdram_s1 => niosII_system_burst_11_downstream_qualified_request_sdram_s1,
      niosII_system_burst_11_downstream_read_data_valid_sdram_s1 => niosII_system_burst_11_downstream_read_data_valid_sdram_s1,
      niosII_system_burst_11_downstream_read_data_valid_sdram_s1_shift_register => niosII_system_burst_11_downstream_read_data_valid_sdram_s1_shift_register,
      niosII_system_burst_11_downstream_requests_sdram_s1 => niosII_system_burst_11_downstream_requests_sdram_s1,
      sdram_s1_address => sdram_s1_address,
      sdram_s1_byteenable_n => sdram_s1_byteenable_n,
      sdram_s1_chipselect => sdram_s1_chipselect,
      sdram_s1_read_n => sdram_s1_read_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_reset_n => sdram_s1_reset_n,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa,
      sdram_s1_write_n => sdram_s1_write_n,
      sdram_s1_writedata => sdram_s1_writedata,
      clk => internal_altpll_inst_c1_out,
      niosII_system_burst_10_downstream_address_to_slave => niosII_system_burst_10_downstream_address_to_slave,
      niosII_system_burst_10_downstream_arbitrationshare => niosII_system_burst_10_downstream_arbitrationshare,
      niosII_system_burst_10_downstream_burstcount => niosII_system_burst_10_downstream_burstcount,
      niosII_system_burst_10_downstream_byteenable => niosII_system_burst_10_downstream_byteenable,
      niosII_system_burst_10_downstream_latency_counter => niosII_system_burst_10_downstream_latency_counter,
      niosII_system_burst_10_downstream_read => niosII_system_burst_10_downstream_read,
      niosII_system_burst_10_downstream_write => niosII_system_burst_10_downstream_write,
      niosII_system_burst_10_downstream_writedata => niosII_system_burst_10_downstream_writedata,
      niosII_system_burst_11_downstream_address_to_slave => niosII_system_burst_11_downstream_address_to_slave,
      niosII_system_burst_11_downstream_arbitrationshare => niosII_system_burst_11_downstream_arbitrationshare,
      niosII_system_burst_11_downstream_burstcount => niosII_system_burst_11_downstream_burstcount,
      niosII_system_burst_11_downstream_byteenable => niosII_system_burst_11_downstream_byteenable,
      niosII_system_burst_11_downstream_latency_counter => niosII_system_burst_11_downstream_latency_counter,
      niosII_system_burst_11_downstream_read => niosII_system_burst_11_downstream_read,
      niosII_system_burst_11_downstream_write => niosII_system_burst_11_downstream_write,
      niosII_system_burst_11_downstream_writedata => niosII_system_burst_11_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      sdram_s1_readdata => sdram_s1_readdata,
      sdram_s1_readdatavalid => sdram_s1_readdatavalid,
      sdram_s1_waitrequest => sdram_s1_waitrequest
    );


  --the_sdram, which is an e_ptf_instance
  the_sdram : sdram
    port map(
      za_data => sdram_s1_readdata,
      za_valid => sdram_s1_readdatavalid,
      za_waitrequest => sdram_s1_waitrequest,
      zs_addr => internal_zs_addr_from_the_sdram,
      zs_ba => internal_zs_ba_from_the_sdram,
      zs_cas_n => internal_zs_cas_n_from_the_sdram,
      zs_cke => internal_zs_cke_from_the_sdram,
      zs_cs_n => internal_zs_cs_n_from_the_sdram,
      zs_dq => zs_dq_to_and_from_the_sdram,
      zs_dqm => internal_zs_dqm_from_the_sdram,
      zs_ras_n => internal_zs_ras_n_from_the_sdram,
      zs_we_n => internal_zs_we_n_from_the_sdram,
      az_addr => sdram_s1_address,
      az_be_n => sdram_s1_byteenable_n,
      az_cs => sdram_s1_chipselect,
      az_data => sdram_s1_writedata,
      az_rd_n => sdram_s1_read_n,
      az_wr_n => sdram_s1_write_n,
      clk => internal_altpll_inst_c1_out,
      reset_n => sdram_s1_reset_n
    );


  --the_seven_seg_pio_s1, which is an e_instance
  the_seven_seg_pio_s1 : seven_seg_pio_s1_arbitrator
    port map(
      d1_seven_seg_pio_s1_end_xfer => d1_seven_seg_pio_s1_end_xfer,
      niosII_system_burst_14_downstream_granted_seven_seg_pio_s1 => niosII_system_burst_14_downstream_granted_seven_seg_pio_s1,
      niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1 => niosII_system_burst_14_downstream_qualified_request_seven_seg_pio_s1,
      niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1 => niosII_system_burst_14_downstream_read_data_valid_seven_seg_pio_s1,
      niosII_system_burst_14_downstream_requests_seven_seg_pio_s1 => niosII_system_burst_14_downstream_requests_seven_seg_pio_s1,
      seven_seg_pio_s1_address => seven_seg_pio_s1_address,
      seven_seg_pio_s1_chipselect => seven_seg_pio_s1_chipselect,
      seven_seg_pio_s1_readdata_from_sa => seven_seg_pio_s1_readdata_from_sa,
      seven_seg_pio_s1_reset_n => seven_seg_pio_s1_reset_n,
      seven_seg_pio_s1_write_n => seven_seg_pio_s1_write_n,
      seven_seg_pio_s1_writedata => seven_seg_pio_s1_writedata,
      clk => internal_altpll_inst_c1_out,
      niosII_system_burst_14_downstream_address_to_slave => niosII_system_burst_14_downstream_address_to_slave,
      niosII_system_burst_14_downstream_arbitrationshare => niosII_system_burst_14_downstream_arbitrationshare,
      niosII_system_burst_14_downstream_burstcount => niosII_system_burst_14_downstream_burstcount,
      niosII_system_burst_14_downstream_latency_counter => niosII_system_burst_14_downstream_latency_counter,
      niosII_system_burst_14_downstream_nativeaddress => niosII_system_burst_14_downstream_nativeaddress,
      niosII_system_burst_14_downstream_read => niosII_system_burst_14_downstream_read,
      niosII_system_burst_14_downstream_write => niosII_system_burst_14_downstream_write,
      niosII_system_burst_14_downstream_writedata => niosII_system_burst_14_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      seven_seg_pio_s1_readdata => seven_seg_pio_s1_readdata
    );


  --the_seven_seg_pio, which is an e_ptf_instance
  the_seven_seg_pio : seven_seg_pio
    port map(
      out_port => internal_out_port_from_the_seven_seg_pio,
      readdata => seven_seg_pio_s1_readdata,
      address => seven_seg_pio_s1_address,
      chipselect => seven_seg_pio_s1_chipselect,
      clk => internal_altpll_inst_c1_out,
      reset_n => seven_seg_pio_s1_reset_n,
      write_n => seven_seg_pio_s1_write_n,
      writedata => seven_seg_pio_s1_writedata
    );


  --the_sram_IF_0, which is an e_ptf_instance
  the_sram_IF_0 : sram_IF_0
    port map(
      ats_tsb_data => sram_IF_0_tsb_data,
      coe_sram_address => internal_coe_sram_address_from_the_sram_IF_0,
      coe_sram_chipenable_n => internal_coe_sram_chipenable_n_from_the_sram_IF_0,
      coe_sram_lowerbyte_n => internal_coe_sram_lowerbyte_n_from_the_sram_IF_0,
      coe_sram_outputenable_n => internal_coe_sram_outputenable_n_from_the_sram_IF_0,
      coe_sram_upperbyte_n => internal_coe_sram_upperbyte_n_from_the_sram_IF_0,
      coe_sram_writeenable_n => internal_coe_sram_writeenable_n_from_the_sram_IF_0,
      ats_tsb_address => sram_IF_0_tsb_address (17 DOWNTO 0),
      ats_tsb_byteenable_n => sram_IF_0_tsb_byteenable_n,
      ats_tsb_chipselect_n => sram_IF_0_tsb_chipselect_n,
      ats_tsb_outputenable_n => sram_IF_0_tsb_outputenable_n,
      ats_tsb_write_n => sram_IF_0_tsb_write_n
    );


  --the_switch_s1, which is an e_instance
  the_switch_s1 : switch_s1_arbitrator
    port map(
      d1_switch_s1_end_xfer => d1_switch_s1_end_xfer,
      niosII_system_burst_9_downstream_granted_switch_s1 => niosII_system_burst_9_downstream_granted_switch_s1,
      niosII_system_burst_9_downstream_qualified_request_switch_s1 => niosII_system_burst_9_downstream_qualified_request_switch_s1,
      niosII_system_burst_9_downstream_read_data_valid_switch_s1 => niosII_system_burst_9_downstream_read_data_valid_switch_s1,
      niosII_system_burst_9_downstream_requests_switch_s1 => niosII_system_burst_9_downstream_requests_switch_s1,
      switch_s1_address => switch_s1_address,
      switch_s1_readdata_from_sa => switch_s1_readdata_from_sa,
      switch_s1_reset_n => switch_s1_reset_n,
      clk => internal_altpll_inst_c1_out,
      niosII_system_burst_9_downstream_address_to_slave => niosII_system_burst_9_downstream_address_to_slave,
      niosII_system_burst_9_downstream_arbitrationshare => niosII_system_burst_9_downstream_arbitrationshare,
      niosII_system_burst_9_downstream_burstcount => niosII_system_burst_9_downstream_burstcount,
      niosII_system_burst_9_downstream_latency_counter => niosII_system_burst_9_downstream_latency_counter,
      niosII_system_burst_9_downstream_nativeaddress => niosII_system_burst_9_downstream_nativeaddress,
      niosII_system_burst_9_downstream_read => niosII_system_burst_9_downstream_read,
      niosII_system_burst_9_downstream_write => niosII_system_burst_9_downstream_write,
      reset_n => altpll_inst_c1_out_reset_n,
      switch_s1_readdata => switch_s1_readdata
    );


  --the_switch, which is an e_ptf_instance
  the_switch : switch
    port map(
      readdata => switch_s1_readdata,
      address => switch_s1_address,
      clk => internal_altpll_inst_c1_out,
      in_port => in_port_to_the_switch,
      reset_n => switch_s1_reset_n
    );


  --the_sys_clk_timer_s1, which is an e_instance
  the_sys_clk_timer_s1 : sys_clk_timer_s1_arbitrator
    port map(
      d1_sys_clk_timer_s1_end_xfer => d1_sys_clk_timer_s1_end_xfer,
      niosII_system_burst_5_downstream_granted_sys_clk_timer_s1 => niosII_system_burst_5_downstream_granted_sys_clk_timer_s1,
      niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1 => niosII_system_burst_5_downstream_qualified_request_sys_clk_timer_s1,
      niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1 => niosII_system_burst_5_downstream_read_data_valid_sys_clk_timer_s1,
      niosII_system_burst_5_downstream_requests_sys_clk_timer_s1 => niosII_system_burst_5_downstream_requests_sys_clk_timer_s1,
      sys_clk_timer_s1_address => sys_clk_timer_s1_address,
      sys_clk_timer_s1_chipselect => sys_clk_timer_s1_chipselect,
      sys_clk_timer_s1_irq_from_sa => sys_clk_timer_s1_irq_from_sa,
      sys_clk_timer_s1_readdata_from_sa => sys_clk_timer_s1_readdata_from_sa,
      sys_clk_timer_s1_reset_n => sys_clk_timer_s1_reset_n,
      sys_clk_timer_s1_write_n => sys_clk_timer_s1_write_n,
      sys_clk_timer_s1_writedata => sys_clk_timer_s1_writedata,
      clk => internal_altpll_inst_c1_out,
      niosII_system_burst_5_downstream_address_to_slave => niosII_system_burst_5_downstream_address_to_slave,
      niosII_system_burst_5_downstream_arbitrationshare => niosII_system_burst_5_downstream_arbitrationshare,
      niosII_system_burst_5_downstream_burstcount => niosII_system_burst_5_downstream_burstcount,
      niosII_system_burst_5_downstream_latency_counter => niosII_system_burst_5_downstream_latency_counter,
      niosII_system_burst_5_downstream_nativeaddress => niosII_system_burst_5_downstream_nativeaddress,
      niosII_system_burst_5_downstream_read => niosII_system_burst_5_downstream_read,
      niosII_system_burst_5_downstream_write => niosII_system_burst_5_downstream_write,
      niosII_system_burst_5_downstream_writedata => niosII_system_burst_5_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      sys_clk_timer_s1_irq => sys_clk_timer_s1_irq,
      sys_clk_timer_s1_readdata => sys_clk_timer_s1_readdata
    );


  --the_sys_clk_timer, which is an e_ptf_instance
  the_sys_clk_timer : sys_clk_timer
    port map(
      irq => sys_clk_timer_s1_irq,
      readdata => sys_clk_timer_s1_readdata,
      address => sys_clk_timer_s1_address,
      chipselect => sys_clk_timer_s1_chipselect,
      clk => internal_altpll_inst_c1_out,
      reset_n => sys_clk_timer_s1_reset_n,
      write_n => sys_clk_timer_s1_write_n,
      writedata => sys_clk_timer_s1_writedata
    );


  --the_sysid_control_slave, which is an e_instance
  the_sysid_control_slave : sysid_control_slave_arbitrator
    port map(
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      niosII_system_burst_4_downstream_granted_sysid_control_slave => niosII_system_burst_4_downstream_granted_sysid_control_slave,
      niosII_system_burst_4_downstream_qualified_request_sysid_control_slave => niosII_system_burst_4_downstream_qualified_request_sysid_control_slave,
      niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave => niosII_system_burst_4_downstream_read_data_valid_sysid_control_slave,
      niosII_system_burst_4_downstream_requests_sysid_control_slave => niosII_system_burst_4_downstream_requests_sysid_control_slave,
      sysid_control_slave_address => sysid_control_slave_address,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa,
      sysid_control_slave_reset_n => sysid_control_slave_reset_n,
      clk => internal_altpll_inst_c1_out,
      niosII_system_burst_4_downstream_address_to_slave => niosII_system_burst_4_downstream_address_to_slave,
      niosII_system_burst_4_downstream_arbitrationshare => niosII_system_burst_4_downstream_arbitrationshare,
      niosII_system_burst_4_downstream_burstcount => niosII_system_burst_4_downstream_burstcount,
      niosII_system_burst_4_downstream_latency_counter => niosII_system_burst_4_downstream_latency_counter,
      niosII_system_burst_4_downstream_nativeaddress => niosII_system_burst_4_downstream_nativeaddress,
      niosII_system_burst_4_downstream_read => niosII_system_burst_4_downstream_read,
      niosII_system_burst_4_downstream_write => niosII_system_burst_4_downstream_write,
      reset_n => altpll_inst_c1_out_reset_n,
      sysid_control_slave_readdata => sysid_control_slave_readdata
    );


  --the_sysid, which is an e_ptf_instance
  the_sysid : sysid
    port map(
      readdata => sysid_control_slave_readdata,
      address => sysid_control_slave_address,
      clock => sysid_control_slave_clock,
      reset_n => sysid_control_slave_reset_n
    );


  --the_tri_state_bridge_avalon_slave, which is an e_instance
  the_tri_state_bridge_avalon_slave : tri_state_bridge_avalon_slave_arbitrator
    port map(
      address_to_the_ext_flash => internal_address_to_the_ext_flash,
      d1_tri_state_bridge_avalon_slave_end_xfer => d1_tri_state_bridge_avalon_slave_end_xfer,
      data_to_and_from_the_ext_flash => data_to_and_from_the_ext_flash,
      ext_flash_s1_wait_counter_eq_0 => ext_flash_s1_wait_counter_eq_0,
      incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0 => incoming_data_to_and_from_the_ext_flash_with_Xs_converted_to_0,
      niosII_system_burst_12_downstream_granted_ext_flash_s1 => niosII_system_burst_12_downstream_granted_ext_flash_s1,
      niosII_system_burst_12_downstream_qualified_request_ext_flash_s1 => niosII_system_burst_12_downstream_qualified_request_ext_flash_s1,
      niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1 => niosII_system_burst_12_downstream_read_data_valid_ext_flash_s1,
      niosII_system_burst_12_downstream_requests_ext_flash_s1 => niosII_system_burst_12_downstream_requests_ext_flash_s1,
      niosII_system_burst_13_downstream_granted_ext_flash_s1 => niosII_system_burst_13_downstream_granted_ext_flash_s1,
      niosII_system_burst_13_downstream_qualified_request_ext_flash_s1 => niosII_system_burst_13_downstream_qualified_request_ext_flash_s1,
      niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1 => niosII_system_burst_13_downstream_read_data_valid_ext_flash_s1,
      niosII_system_burst_13_downstream_requests_ext_flash_s1 => niosII_system_burst_13_downstream_requests_ext_flash_s1,
      read_n_to_the_ext_flash => internal_read_n_to_the_ext_flash,
      select_n_to_the_ext_flash => internal_select_n_to_the_ext_flash,
      write_n_to_the_ext_flash => internal_write_n_to_the_ext_flash,
      clk => internal_altpll_inst_c1_out,
      niosII_system_burst_12_downstream_address_to_slave => niosII_system_burst_12_downstream_address_to_slave,
      niosII_system_burst_12_downstream_arbitrationshare => niosII_system_burst_12_downstream_arbitrationshare,
      niosII_system_burst_12_downstream_burstcount => niosII_system_burst_12_downstream_burstcount,
      niosII_system_burst_12_downstream_byteenable => niosII_system_burst_12_downstream_byteenable,
      niosII_system_burst_12_downstream_latency_counter => niosII_system_burst_12_downstream_latency_counter,
      niosII_system_burst_12_downstream_read => niosII_system_burst_12_downstream_read,
      niosII_system_burst_12_downstream_write => niosII_system_burst_12_downstream_write,
      niosII_system_burst_12_downstream_writedata => niosII_system_burst_12_downstream_writedata,
      niosII_system_burst_13_downstream_address_to_slave => niosII_system_burst_13_downstream_address_to_slave,
      niosII_system_burst_13_downstream_arbitrationshare => niosII_system_burst_13_downstream_arbitrationshare,
      niosII_system_burst_13_downstream_burstcount => niosII_system_burst_13_downstream_burstcount,
      niosII_system_burst_13_downstream_byteenable => niosII_system_burst_13_downstream_byteenable,
      niosII_system_burst_13_downstream_latency_counter => niosII_system_burst_13_downstream_latency_counter,
      niosII_system_burst_13_downstream_read => niosII_system_burst_13_downstream_read,
      niosII_system_burst_13_downstream_write => niosII_system_burst_13_downstream_write,
      niosII_system_burst_13_downstream_writedata => niosII_system_burst_13_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_tsb_avalon_slave, which is an e_instance
  the_tsb_avalon_slave : tsb_avalon_slave_arbitrator
    port map(
      d1_tsb_avalon_slave_end_xfer => d1_tsb_avalon_slave_end_xfer,
      incoming_sram_IF_0_tsb_data => incoming_sram_IF_0_tsb_data,
      niosII_system_burst_19_downstream_granted_sram_IF_0_tsb => niosII_system_burst_19_downstream_granted_sram_IF_0_tsb,
      niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb => niosII_system_burst_19_downstream_qualified_request_sram_IF_0_tsb,
      niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb => niosII_system_burst_19_downstream_read_data_valid_sram_IF_0_tsb,
      niosII_system_burst_19_downstream_requests_sram_IF_0_tsb => niosII_system_burst_19_downstream_requests_sram_IF_0_tsb,
      niosII_system_burst_20_downstream_granted_sram_IF_0_tsb => niosII_system_burst_20_downstream_granted_sram_IF_0_tsb,
      niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb => niosII_system_burst_20_downstream_qualified_request_sram_IF_0_tsb,
      niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb => niosII_system_burst_20_downstream_read_data_valid_sram_IF_0_tsb,
      niosII_system_burst_20_downstream_requests_sram_IF_0_tsb => niosII_system_burst_20_downstream_requests_sram_IF_0_tsb,
      sram_IF_0_tsb_address => sram_IF_0_tsb_address,
      sram_IF_0_tsb_byteenable_n => sram_IF_0_tsb_byteenable_n,
      sram_IF_0_tsb_chipselect_n => sram_IF_0_tsb_chipselect_n,
      sram_IF_0_tsb_data => sram_IF_0_tsb_data,
      sram_IF_0_tsb_outputenable_n => sram_IF_0_tsb_outputenable_n,
      sram_IF_0_tsb_write_n => sram_IF_0_tsb_write_n,
      clk => internal_altpll_inst_c1_out,
      niosII_system_burst_19_downstream_address_to_slave => niosII_system_burst_19_downstream_address_to_slave,
      niosII_system_burst_19_downstream_arbitrationshare => niosII_system_burst_19_downstream_arbitrationshare,
      niosII_system_burst_19_downstream_burstcount => niosII_system_burst_19_downstream_burstcount,
      niosII_system_burst_19_downstream_byteenable => niosII_system_burst_19_downstream_byteenable,
      niosII_system_burst_19_downstream_latency_counter => niosII_system_burst_19_downstream_latency_counter,
      niosII_system_burst_19_downstream_read => niosII_system_burst_19_downstream_read,
      niosII_system_burst_19_downstream_write => niosII_system_burst_19_downstream_write,
      niosII_system_burst_19_downstream_writedata => niosII_system_burst_19_downstream_writedata,
      niosII_system_burst_20_downstream_address_to_slave => niosII_system_burst_20_downstream_address_to_slave,
      niosII_system_burst_20_downstream_arbitrationshare => niosII_system_burst_20_downstream_arbitrationshare,
      niosII_system_burst_20_downstream_burstcount => niosII_system_burst_20_downstream_burstcount,
      niosII_system_burst_20_downstream_byteenable => niosII_system_burst_20_downstream_byteenable,
      niosII_system_burst_20_downstream_latency_counter => niosII_system_burst_20_downstream_latency_counter,
      niosII_system_burst_20_downstream_read => niosII_system_burst_20_downstream_read,
      niosII_system_burst_20_downstream_write => niosII_system_burst_20_downstream_write,
      niosII_system_burst_20_downstream_writedata => niosII_system_burst_20_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n
    );


  --the_uart_0_s1, which is an e_instance
  the_uart_0_s1 : uart_0_s1_arbitrator
    port map(
      d1_uart_0_s1_end_xfer => d1_uart_0_s1_end_xfer,
      niosII_system_burst_17_downstream_granted_uart_0_s1 => niosII_system_burst_17_downstream_granted_uart_0_s1,
      niosII_system_burst_17_downstream_qualified_request_uart_0_s1 => niosII_system_burst_17_downstream_qualified_request_uart_0_s1,
      niosII_system_burst_17_downstream_read_data_valid_uart_0_s1 => niosII_system_burst_17_downstream_read_data_valid_uart_0_s1,
      niosII_system_burst_17_downstream_requests_uart_0_s1 => niosII_system_burst_17_downstream_requests_uart_0_s1,
      uart_0_s1_address => uart_0_s1_address,
      uart_0_s1_begintransfer => uart_0_s1_begintransfer,
      uart_0_s1_chipselect => uart_0_s1_chipselect,
      uart_0_s1_dataavailable_from_sa => uart_0_s1_dataavailable_from_sa,
      uart_0_s1_irq_from_sa => uart_0_s1_irq_from_sa,
      uart_0_s1_read_n => uart_0_s1_read_n,
      uart_0_s1_readdata_from_sa => uart_0_s1_readdata_from_sa,
      uart_0_s1_readyfordata_from_sa => uart_0_s1_readyfordata_from_sa,
      uart_0_s1_reset_n => uart_0_s1_reset_n,
      uart_0_s1_write_n => uart_0_s1_write_n,
      uart_0_s1_writedata => uart_0_s1_writedata,
      clk => internal_altpll_inst_c1_out,
      niosII_system_burst_17_downstream_address_to_slave => niosII_system_burst_17_downstream_address_to_slave,
      niosII_system_burst_17_downstream_arbitrationshare => niosII_system_burst_17_downstream_arbitrationshare,
      niosII_system_burst_17_downstream_burstcount => niosII_system_burst_17_downstream_burstcount,
      niosII_system_burst_17_downstream_latency_counter => niosII_system_burst_17_downstream_latency_counter,
      niosII_system_burst_17_downstream_nativeaddress => niosII_system_burst_17_downstream_nativeaddress,
      niosII_system_burst_17_downstream_read => niosII_system_burst_17_downstream_read,
      niosII_system_burst_17_downstream_write => niosII_system_burst_17_downstream_write,
      niosII_system_burst_17_downstream_writedata => niosII_system_burst_17_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      uart_0_s1_dataavailable => uart_0_s1_dataavailable,
      uart_0_s1_irq => uart_0_s1_irq,
      uart_0_s1_readdata => uart_0_s1_readdata,
      uart_0_s1_readyfordata => uart_0_s1_readyfordata
    );


  --the_uart_0, which is an e_ptf_instance
  the_uart_0 : uart_0
    port map(
      dataavailable => uart_0_s1_dataavailable,
      irq => uart_0_s1_irq,
      readdata => uart_0_s1_readdata,
      readyfordata => uart_0_s1_readyfordata,
      txd => internal_txd_from_the_uart_0,
      address => uart_0_s1_address,
      begintransfer => uart_0_s1_begintransfer,
      chipselect => uart_0_s1_chipselect,
      clk => internal_altpll_inst_c1_out,
      read_n => uart_0_s1_read_n,
      reset_n => uart_0_s1_reset_n,
      rxd => rxd_to_the_uart_0,
      write_n => uart_0_s1_write_n,
      writedata => uart_0_s1_writedata
    );


  --the_uart_1_s1, which is an e_instance
  the_uart_1_s1 : uart_1_s1_arbitrator
    port map(
      d1_uart_1_s1_end_xfer => d1_uart_1_s1_end_xfer,
      niosII_system_burst_18_downstream_granted_uart_1_s1 => niosII_system_burst_18_downstream_granted_uart_1_s1,
      niosII_system_burst_18_downstream_qualified_request_uart_1_s1 => niosII_system_burst_18_downstream_qualified_request_uart_1_s1,
      niosII_system_burst_18_downstream_read_data_valid_uart_1_s1 => niosII_system_burst_18_downstream_read_data_valid_uart_1_s1,
      niosII_system_burst_18_downstream_requests_uart_1_s1 => niosII_system_burst_18_downstream_requests_uart_1_s1,
      uart_1_s1_address => uart_1_s1_address,
      uart_1_s1_begintransfer => uart_1_s1_begintransfer,
      uart_1_s1_chipselect => uart_1_s1_chipselect,
      uart_1_s1_dataavailable_from_sa => uart_1_s1_dataavailable_from_sa,
      uart_1_s1_irq_from_sa => uart_1_s1_irq_from_sa,
      uart_1_s1_read_n => uart_1_s1_read_n,
      uart_1_s1_readdata_from_sa => uart_1_s1_readdata_from_sa,
      uart_1_s1_readyfordata_from_sa => uart_1_s1_readyfordata_from_sa,
      uart_1_s1_reset_n => uart_1_s1_reset_n,
      uart_1_s1_write_n => uart_1_s1_write_n,
      uart_1_s1_writedata => uart_1_s1_writedata,
      clk => internal_altpll_inst_c1_out,
      niosII_system_burst_18_downstream_address_to_slave => niosII_system_burst_18_downstream_address_to_slave,
      niosII_system_burst_18_downstream_arbitrationshare => niosII_system_burst_18_downstream_arbitrationshare,
      niosII_system_burst_18_downstream_burstcount => niosII_system_burst_18_downstream_burstcount,
      niosII_system_burst_18_downstream_latency_counter => niosII_system_burst_18_downstream_latency_counter,
      niosII_system_burst_18_downstream_nativeaddress => niosII_system_burst_18_downstream_nativeaddress,
      niosII_system_burst_18_downstream_read => niosII_system_burst_18_downstream_read,
      niosII_system_burst_18_downstream_write => niosII_system_burst_18_downstream_write,
      niosII_system_burst_18_downstream_writedata => niosII_system_burst_18_downstream_writedata,
      reset_n => altpll_inst_c1_out_reset_n,
      uart_1_s1_dataavailable => uart_1_s1_dataavailable,
      uart_1_s1_irq => uart_1_s1_irq,
      uart_1_s1_readdata => uart_1_s1_readdata,
      uart_1_s1_readyfordata => uart_1_s1_readyfordata
    );


  --the_uart_1, which is an e_ptf_instance
  the_uart_1 : uart_1
    port map(
      dataavailable => uart_1_s1_dataavailable,
      irq => uart_1_s1_irq,
      readdata => uart_1_s1_readdata,
      readyfordata => uart_1_s1_readyfordata,
      txd => internal_txd_from_the_uart_1,
      address => uart_1_s1_address,
      begintransfer => uart_1_s1_begintransfer,
      chipselect => uart_1_s1_chipselect,
      clk => internal_altpll_inst_c1_out,
      read_n => uart_1_s1_read_n,
      reset_n => uart_1_s1_reset_n,
      rxd => rxd_to_the_uart_1,
      write_n => uart_1_s1_write_n,
      writedata => uart_1_s1_writedata
    );


  --reset is asserted asynchronously and deasserted synchronously
  niosII_system_reset_clk_0_domain_synch : niosII_system_reset_clk_0_domain_synch_module
    port map(
      data_out => clk_0_reset_n,
      clk => clk_0,
      data_in => module_input138,
      reset_n => reset_n_sources
    );

  module_input138 <= std_logic'('1');

  --reset sources mux, which is an e_mux
  reset_n_sources <= Vector_To_Std_Logic(NOT ((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT reset_n))) OR std_logic_vector'("00000000000000000000000000000000")) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_resetrequest_from_sa))))));
  --reset is asserted asynchronously and deasserted synchronously
  niosII_system_reset_altpll_inst_c1_out_domain_synch : niosII_system_reset_altpll_inst_c1_out_domain_synch_module
    port map(
      data_out => altpll_inst_c1_out_reset_n,
      clk => internal_altpll_inst_c1_out,
      data_in => module_input139,
      reset_n => reset_n_sources
    );

  module_input139 <= std_logic'('1');

  --niosII_system_burst_0_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  niosII_system_burst_0_upstream_writedata <= std_logic_vector'("00000000000000000000000000000000");
  --niosII_system_burst_10_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  niosII_system_burst_10_upstream_writedata <= std_logic_vector'("0000000000000000");
  --niosII_system_burst_12_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  niosII_system_burst_12_upstream_writedata <= std_logic_vector'("00000000");
  --niosII_system_burst_19_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  niosII_system_burst_19_upstream_writedata <= std_logic_vector'("0000000000000000");
  --niosII_system_burst_2_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  niosII_system_burst_2_upstream_writedata <= std_logic_vector'("00000000000000000000000000000000");
  --niosII_system_clock_0_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  niosII_system_clock_0_out_endofpacket <= std_logic'('0');
  --sysid_control_slave_clock of type clock does not connect to anything so wire it to default (0)
  sysid_control_slave_clock <= std_logic'('0');
  --vhdl renameroo for output signals
  ENET_CMD_from_the_dm9000a_inst <= internal_ENET_CMD_from_the_dm9000a_inst;
  --vhdl renameroo for output signals
  ENET_CS_N_from_the_dm9000a_inst <= internal_ENET_CS_N_from_the_dm9000a_inst;
  --vhdl renameroo for output signals
  ENET_RD_N_from_the_dm9000a_inst <= internal_ENET_RD_N_from_the_dm9000a_inst;
  --vhdl renameroo for output signals
  ENET_RST_N_from_the_dm9000a_inst <= internal_ENET_RST_N_from_the_dm9000a_inst;
  --vhdl renameroo for output signals
  ENET_WR_N_from_the_dm9000a_inst <= internal_ENET_WR_N_from_the_dm9000a_inst;
  --vhdl renameroo for output signals
  LCD_E_from_the_lcd_display <= internal_LCD_E_from_the_lcd_display;
  --vhdl renameroo for output signals
  LCD_RS_from_the_lcd_display <= internal_LCD_RS_from_the_lcd_display;
  --vhdl renameroo for output signals
  LCD_RW_from_the_lcd_display <= internal_LCD_RW_from_the_lcd_display;
  --vhdl renameroo for output signals
  address_to_the_ext_flash <= internal_address_to_the_ext_flash;
  --vhdl renameroo for output signals
  altpll_inst_c1_out <= internal_altpll_inst_c1_out;
  --vhdl renameroo for output signals
  coe_sram_address_from_the_sram_IF_0 <= internal_coe_sram_address_from_the_sram_IF_0;
  --vhdl renameroo for output signals
  coe_sram_chipenable_n_from_the_sram_IF_0 <= internal_coe_sram_chipenable_n_from_the_sram_IF_0;
  --vhdl renameroo for output signals
  coe_sram_lowerbyte_n_from_the_sram_IF_0 <= internal_coe_sram_lowerbyte_n_from_the_sram_IF_0;
  --vhdl renameroo for output signals
  coe_sram_outputenable_n_from_the_sram_IF_0 <= internal_coe_sram_outputenable_n_from_the_sram_IF_0;
  --vhdl renameroo for output signals
  coe_sram_upperbyte_n_from_the_sram_IF_0 <= internal_coe_sram_upperbyte_n_from_the_sram_IF_0;
  --vhdl renameroo for output signals
  coe_sram_writeenable_n_from_the_sram_IF_0 <= internal_coe_sram_writeenable_n_from_the_sram_IF_0;
  --vhdl renameroo for output signals
  locked_from_the_altpll_inst <= internal_locked_from_the_altpll_inst;
  --vhdl renameroo for output signals
  out_port_from_the_led_pio <= internal_out_port_from_the_led_pio;
  --vhdl renameroo for output signals
  out_port_from_the_seven_seg_pio <= internal_out_port_from_the_seven_seg_pio;
  --vhdl renameroo for output signals
  phasedone_from_the_altpll_inst <= internal_phasedone_from_the_altpll_inst;
  --vhdl renameroo for output signals
  read_n_to_the_ext_flash <= internal_read_n_to_the_ext_flash;
  --vhdl renameroo for output signals
  select_n_to_the_ext_flash <= internal_select_n_to_the_ext_flash;
  --vhdl renameroo for output signals
  txd_from_the_uart_0 <= internal_txd_from_the_uart_0;
  --vhdl renameroo for output signals
  txd_from_the_uart_1 <= internal_txd_from_the_uart_1;
  --vhdl renameroo for output signals
  write_n_to_the_ext_flash <= internal_write_n_to_the_ext_flash;
  --vhdl renameroo for output signals
  zs_addr_from_the_sdram <= internal_zs_addr_from_the_sdram;
  --vhdl renameroo for output signals
  zs_ba_from_the_sdram <= internal_zs_ba_from_the_sdram;
  --vhdl renameroo for output signals
  zs_cas_n_from_the_sdram <= internal_zs_cas_n_from_the_sdram;
  --vhdl renameroo for output signals
  zs_cke_from_the_sdram <= internal_zs_cke_from_the_sdram;
  --vhdl renameroo for output signals
  zs_cs_n_from_the_sdram <= internal_zs_cs_n_from_the_sdram;
  --vhdl renameroo for output signals
  zs_dqm_from_the_sdram <= internal_zs_dqm_from_the_sdram;
  --vhdl renameroo for output signals
  zs_ras_n_from_the_sdram <= internal_zs_ras_n_from_the_sdram;
  --vhdl renameroo for output signals
  zs_we_n_from_the_sdram <= internal_zs_we_n_from_the_sdram;

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ext_flash_lane0_module is 
        port (
              -- inputs:
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ext_flash_lane0_module;


architecture europa of ext_flash_lane0_module is
              signal internal_q :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 4194303 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, rdaddress) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (21 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "ext_flash.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 4194304) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rdaddress)));
      


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity ext_flash_lane0_module is 
--        port (
--              
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity ext_flash_lane0_module;
--
--
--architecture europa of ext_flash_lane0_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal internal_q :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 4194303 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
--
--begin
--
--  process (rdaddress)
--  begin
--      read_address <= rdaddress;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "ext_flash.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "UNREGISTERED",
--      lpm_rdaddress_control => "UNREGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 22,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ext_flash is 
        port (
              -- inputs:
                 signal address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal read_n : IN STD_LOGIC;
                 signal select_n : IN STD_LOGIC;
                 signal write_n : IN STD_LOGIC;

              -- outputs:
                 signal data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ext_flash;


architecture europa of ext_flash is
--synthesis translate_off
component ext_flash_lane0_module is 
           port (
                 -- inputs:
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ext_flash_lane0_module;

--synthesis translate_on
                signal data_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal logic_vector_gasket :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal module_input140 :  STD_LOGIC;
                signal module_input141 :  STD_LOGIC;
                signal q_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);

begin

  --s1, which is an e_ptf_slave
--synthesis translate_off
    logic_vector_gasket <= data;
    data_0 <= logic_vector_gasket(7 DOWNTO 0);
    --ext_flash_lane0, which is an e_ram
    ext_flash_lane0 : ext_flash_lane0_module
      port map(
        q => q_0,
        data => data_0,
        rdaddress => address,
        rdclken => module_input140,
        wraddress => address,
        wrclock => write_n,
        wren => module_input141
      );

    module_input140 <= std_logic'('1');
    module_input141 <= NOT select_n;

    data <= A_WE_StdLogicVector((std_logic'(((NOT select_n AND NOT read_n))) = '1'), q_0, A_REP(std_logic'('Z'), 8));
--synthesis translate_on

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your libraries here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>

entity test_bench is 
end entity test_bench;


architecture europa of test_bench is
component niosII_system is 
           port (
                 -- 1) global signals:
                    signal altpll_inst_c0_out : OUT STD_LOGIC;
                    signal altpll_inst_c1_out : OUT STD_LOGIC;
                    signal altpll_inst_c2_out : OUT STD_LOGIC;
                    signal clk_0 : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sram_IF_0_tsb_data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_altpll_inst
                    signal locked_from_the_altpll_inst : OUT STD_LOGIC;
                    signal phasedone_from_the_altpll_inst : OUT STD_LOGIC;

                 -- the_dm9000a_inst
                    signal ENET_CMD_from_the_dm9000a_inst : OUT STD_LOGIC;
                    signal ENET_CS_N_from_the_dm9000a_inst : OUT STD_LOGIC;
                    signal ENET_DATA_to_and_from_the_dm9000a_inst : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal ENET_INT_to_the_dm9000a_inst : IN STD_LOGIC;
                    signal ENET_RD_N_from_the_dm9000a_inst : OUT STD_LOGIC;
                    signal ENET_RST_N_from_the_dm9000a_inst : OUT STD_LOGIC;
                    signal ENET_WR_N_from_the_dm9000a_inst : OUT STD_LOGIC;

                 -- the_lcd_display
                    signal LCD_E_from_the_lcd_display : OUT STD_LOGIC;
                    signal LCD_RS_from_the_lcd_display : OUT STD_LOGIC;
                    signal LCD_RW_from_the_lcd_display : OUT STD_LOGIC;
                    signal LCD_data_to_and_from_the_lcd_display : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_led_pio
                    signal out_port_from_the_led_pio : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_sdram
                    signal zs_addr_from_the_sdram : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n_from_the_sdram : OUT STD_LOGIC;
                    signal zs_cke_from_the_sdram : OUT STD_LOGIC;
                    signal zs_cs_n_from_the_sdram : OUT STD_LOGIC;
                    signal zs_dq_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal zs_dqm_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n_from_the_sdram : OUT STD_LOGIC;
                    signal zs_we_n_from_the_sdram : OUT STD_LOGIC;

                 -- the_seven_seg_pio
                    signal out_port_from_the_seven_seg_pio : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_sram_IF_0
                    signal coe_sram_address_from_the_sram_IF_0 : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal coe_sram_chipenable_n_from_the_sram_IF_0 : OUT STD_LOGIC;
                    signal coe_sram_lowerbyte_n_from_the_sram_IF_0 : OUT STD_LOGIC;
                    signal coe_sram_outputenable_n_from_the_sram_IF_0 : OUT STD_LOGIC;
                    signal coe_sram_upperbyte_n_from_the_sram_IF_0 : OUT STD_LOGIC;
                    signal coe_sram_writeenable_n_from_the_sram_IF_0 : OUT STD_LOGIC;

                 -- the_switch
                    signal in_port_to_the_switch : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_tri_state_bridge_avalon_slave
                    signal address_to_the_ext_flash : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal data_to_and_from_the_ext_flash : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal read_n_to_the_ext_flash : OUT STD_LOGIC;
                    signal select_n_to_the_ext_flash : OUT STD_LOGIC;
                    signal write_n_to_the_ext_flash : OUT STD_LOGIC;

                 -- the_uart_0
                    signal rxd_to_the_uart_0 : IN STD_LOGIC;
                    signal txd_from_the_uart_0 : OUT STD_LOGIC;

                 -- the_uart_1
                    signal rxd_to_the_uart_1 : IN STD_LOGIC;
                    signal txd_from_the_uart_1 : OUT STD_LOGIC
                 );
end component niosII_system;

component ext_flash is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal read_n : IN STD_LOGIC;
                    signal select_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;

                 -- outputs:
                    signal data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ext_flash;

                signal ENET_CMD_from_the_dm9000a_inst :  STD_LOGIC;
                signal ENET_CS_N_from_the_dm9000a_inst :  STD_LOGIC;
                signal ENET_DATA_to_and_from_the_dm9000a_inst :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal ENET_INT_to_the_dm9000a_inst :  STD_LOGIC;
                signal ENET_RD_N_from_the_dm9000a_inst :  STD_LOGIC;
                signal ENET_RST_N_from_the_dm9000a_inst :  STD_LOGIC;
                signal ENET_WR_N_from_the_dm9000a_inst :  STD_LOGIC;
                signal LCD_E_from_the_lcd_display :  STD_LOGIC;
                signal LCD_RS_from_the_lcd_display :  STD_LOGIC;
                signal LCD_RW_from_the_lcd_display :  STD_LOGIC;
                signal LCD_data_to_and_from_the_lcd_display :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal address_to_the_ext_flash :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal altpll_inst_c0_out :  STD_LOGIC;
                signal altpll_inst_c1_out :  STD_LOGIC;
                signal altpll_inst_c2_out :  STD_LOGIC;
                signal clk :  STD_LOGIC;
                signal clk_0 :  STD_LOGIC;
                signal coe_sram_address_from_the_sram_IF_0 :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal coe_sram_chipenable_n_from_the_sram_IF_0 :  STD_LOGIC;
                signal coe_sram_lowerbyte_n_from_the_sram_IF_0 :  STD_LOGIC;
                signal coe_sram_outputenable_n_from_the_sram_IF_0 :  STD_LOGIC;
                signal coe_sram_upperbyte_n_from_the_sram_IF_0 :  STD_LOGIC;
                signal coe_sram_writeenable_n_from_the_sram_IF_0 :  STD_LOGIC;
                signal data_to_and_from_the_ext_flash :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal in_port_to_the_switch :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal locked_from_the_altpll_inst :  STD_LOGIC;
                signal niosII_system_burst_0_downstream_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_0_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_10_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_10_downstream_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_10_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_11_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_11_downstream_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal niosII_system_burst_12_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_12_downstream_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_12_upstream_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_system_burst_13_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_13_downstream_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal niosII_system_burst_14_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_15_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_16_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_17_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_18_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_19_downstream_nativeaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_19_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_system_burst_1_downstream_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal niosII_system_burst_20_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_20_downstream_nativeaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal niosII_system_burst_21_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_2_downstream_nativeaddress :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_2_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_system_burst_3_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_3_downstream_nativeaddress :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal niosII_system_burst_4_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_5_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_6_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_7_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_8_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_burst_9_downstream_debugaccess :  STD_LOGIC;
                signal niosII_system_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_system_clock_0_out_endofpacket :  STD_LOGIC;
                signal niosII_system_clock_0_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal out_port_from_the_led_pio :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal out_port_from_the_seven_seg_pio :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal phasedone_from_the_altpll_inst :  STD_LOGIC;
                signal read_n_to_the_ext_flash :  STD_LOGIC;
                signal reset_n :  STD_LOGIC;
                signal rxd_to_the_uart_0 :  STD_LOGIC;
                signal rxd_to_the_uart_1 :  STD_LOGIC;
                signal select_n_to_the_ext_flash :  STD_LOGIC;
                signal sram_IF_0_tsb_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sysid_control_slave_clock :  STD_LOGIC;
                signal txd_from_the_uart_0 :  STD_LOGIC;
                signal txd_from_the_uart_1 :  STD_LOGIC;
                signal uart_0_s1_dataavailable_from_sa :  STD_LOGIC;
                signal uart_0_s1_readyfordata_from_sa :  STD_LOGIC;
                signal uart_1_s1_dataavailable_from_sa :  STD_LOGIC;
                signal uart_1_s1_readyfordata_from_sa :  STD_LOGIC;
                signal write_n_to_the_ext_flash :  STD_LOGIC;
                signal zs_addr_from_the_sdram :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal zs_ba_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_cas_n_from_the_sdram :  STD_LOGIC;
                signal zs_cke_from_the_sdram :  STD_LOGIC;
                signal zs_cs_n_from_the_sdram :  STD_LOGIC;
                signal zs_dq_to_and_from_the_sdram :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal zs_dqm_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_ras_n_from_the_sdram :  STD_LOGIC;
                signal zs_we_n_from_the_sdram :  STD_LOGIC;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your component and signal declaration here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


begin

  --Set us up the Dut
  DUT : niosII_system
    port map(
      ENET_CMD_from_the_dm9000a_inst => ENET_CMD_from_the_dm9000a_inst,
      ENET_CS_N_from_the_dm9000a_inst => ENET_CS_N_from_the_dm9000a_inst,
      ENET_DATA_to_and_from_the_dm9000a_inst => ENET_DATA_to_and_from_the_dm9000a_inst,
      ENET_RD_N_from_the_dm9000a_inst => ENET_RD_N_from_the_dm9000a_inst,
      ENET_RST_N_from_the_dm9000a_inst => ENET_RST_N_from_the_dm9000a_inst,
      ENET_WR_N_from_the_dm9000a_inst => ENET_WR_N_from_the_dm9000a_inst,
      LCD_E_from_the_lcd_display => LCD_E_from_the_lcd_display,
      LCD_RS_from_the_lcd_display => LCD_RS_from_the_lcd_display,
      LCD_RW_from_the_lcd_display => LCD_RW_from_the_lcd_display,
      LCD_data_to_and_from_the_lcd_display => LCD_data_to_and_from_the_lcd_display,
      address_to_the_ext_flash => address_to_the_ext_flash,
      altpll_inst_c0_out => altpll_inst_c0_out,
      altpll_inst_c1_out => altpll_inst_c1_out,
      altpll_inst_c2_out => altpll_inst_c2_out,
      coe_sram_address_from_the_sram_IF_0 => coe_sram_address_from_the_sram_IF_0,
      coe_sram_chipenable_n_from_the_sram_IF_0 => coe_sram_chipenable_n_from_the_sram_IF_0,
      coe_sram_lowerbyte_n_from_the_sram_IF_0 => coe_sram_lowerbyte_n_from_the_sram_IF_0,
      coe_sram_outputenable_n_from_the_sram_IF_0 => coe_sram_outputenable_n_from_the_sram_IF_0,
      coe_sram_upperbyte_n_from_the_sram_IF_0 => coe_sram_upperbyte_n_from_the_sram_IF_0,
      coe_sram_writeenable_n_from_the_sram_IF_0 => coe_sram_writeenable_n_from_the_sram_IF_0,
      data_to_and_from_the_ext_flash => data_to_and_from_the_ext_flash,
      locked_from_the_altpll_inst => locked_from_the_altpll_inst,
      out_port_from_the_led_pio => out_port_from_the_led_pio,
      out_port_from_the_seven_seg_pio => out_port_from_the_seven_seg_pio,
      phasedone_from_the_altpll_inst => phasedone_from_the_altpll_inst,
      read_n_to_the_ext_flash => read_n_to_the_ext_flash,
      select_n_to_the_ext_flash => select_n_to_the_ext_flash,
      sram_IF_0_tsb_data => sram_IF_0_tsb_data,
      txd_from_the_uart_0 => txd_from_the_uart_0,
      txd_from_the_uart_1 => txd_from_the_uart_1,
      write_n_to_the_ext_flash => write_n_to_the_ext_flash,
      zs_addr_from_the_sdram => zs_addr_from_the_sdram,
      zs_ba_from_the_sdram => zs_ba_from_the_sdram,
      zs_cas_n_from_the_sdram => zs_cas_n_from_the_sdram,
      zs_cke_from_the_sdram => zs_cke_from_the_sdram,
      zs_cs_n_from_the_sdram => zs_cs_n_from_the_sdram,
      zs_dq_to_and_from_the_sdram => zs_dq_to_and_from_the_sdram,
      zs_dqm_from_the_sdram => zs_dqm_from_the_sdram,
      zs_ras_n_from_the_sdram => zs_ras_n_from_the_sdram,
      zs_we_n_from_the_sdram => zs_we_n_from_the_sdram,
      ENET_INT_to_the_dm9000a_inst => ENET_INT_to_the_dm9000a_inst,
      clk_0 => clk_0,
      in_port_to_the_switch => in_port_to_the_switch,
      reset_n => reset_n,
      rxd_to_the_uart_0 => rxd_to_the_uart_0,
      rxd_to_the_uart_1 => rxd_to_the_uart_1
    );


  --the_ext_flash, which is an e_ptf_instance
  the_ext_flash : ext_flash
    port map(
      data => data_to_and_from_the_ext_flash,
      address => address_to_the_ext_flash,
      read_n => read_n_to_the_ext_flash,
      select_n => select_n_to_the_ext_flash,
      write_n => write_n_to_the_ext_flash
    );


  --default value specified in MODULE switch ptf port section
  in_port_to_the_switch <= std_logic_vector'("00000000");
  process
  begin
    clk_0 <= '0';
    loop
       wait for 10 ns;
       clk_0 <= not clk_0;
    end loop;
  end process;
  PROCESS
    BEGIN
       reset_n <= '0';
       wait for 200 ns;
       reset_n <= '1'; 
    WAIT;
  END PROCESS;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add additional architecture here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


end europa;



--synthesis translate_on
