  --Example instantiation for system 'niosII_system'
  niosII_system_inst : niosII_system
    port map(
      ENET_CMD_from_the_dm9000a_inst => ENET_CMD_from_the_dm9000a_inst,
      ENET_CS_N_from_the_dm9000a_inst => ENET_CS_N_from_the_dm9000a_inst,
      ENET_DATA_to_and_from_the_dm9000a_inst => ENET_DATA_to_and_from_the_dm9000a_inst,
      ENET_RD_N_from_the_dm9000a_inst => ENET_RD_N_from_the_dm9000a_inst,
      ENET_RST_N_from_the_dm9000a_inst => ENET_RST_N_from_the_dm9000a_inst,
      ENET_WR_N_from_the_dm9000a_inst => ENET_WR_N_from_the_dm9000a_inst,
      LCD_E_from_the_lcd_display => LCD_E_from_the_lcd_display,
      LCD_RS_from_the_lcd_display => LCD_RS_from_the_lcd_display,
      LCD_RW_from_the_lcd_display => LCD_RW_from_the_lcd_display,
      LCD_data_to_and_from_the_lcd_display => LCD_data_to_and_from_the_lcd_display,
      address_to_the_ext_flash => address_to_the_ext_flash,
      altpll_inst_c0_out => altpll_inst_c0_out,
      altpll_inst_c1_out => altpll_inst_c1_out,
      altpll_inst_c2_out => altpll_inst_c2_out,
      coe_sram_address_from_the_sram_IF_0 => coe_sram_address_from_the_sram_IF_0,
      coe_sram_chipenable_n_from_the_sram_IF_0 => coe_sram_chipenable_n_from_the_sram_IF_0,
      coe_sram_lowerbyte_n_from_the_sram_IF_0 => coe_sram_lowerbyte_n_from_the_sram_IF_0,
      coe_sram_outputenable_n_from_the_sram_IF_0 => coe_sram_outputenable_n_from_the_sram_IF_0,
      coe_sram_upperbyte_n_from_the_sram_IF_0 => coe_sram_upperbyte_n_from_the_sram_IF_0,
      coe_sram_writeenable_n_from_the_sram_IF_0 => coe_sram_writeenable_n_from_the_sram_IF_0,
      data_to_and_from_the_ext_flash => data_to_and_from_the_ext_flash,
      locked_from_the_altpll_inst => locked_from_the_altpll_inst,
      out_port_from_the_led_pio => out_port_from_the_led_pio,
      out_port_from_the_seven_seg_pio => out_port_from_the_seven_seg_pio,
      phasedone_from_the_altpll_inst => phasedone_from_the_altpll_inst,
      read_n_to_the_ext_flash => read_n_to_the_ext_flash,
      select_n_to_the_ext_flash => select_n_to_the_ext_flash,
      sram_IF_0_tsb_data => sram_IF_0_tsb_data,
      txd_from_the_uart_0 => txd_from_the_uart_0,
      txd_from_the_uart_1 => txd_from_the_uart_1,
      write_n_to_the_ext_flash => write_n_to_the_ext_flash,
      zs_addr_from_the_sdram => zs_addr_from_the_sdram,
      zs_ba_from_the_sdram => zs_ba_from_the_sdram,
      zs_cas_n_from_the_sdram => zs_cas_n_from_the_sdram,
      zs_cke_from_the_sdram => zs_cke_from_the_sdram,
      zs_cs_n_from_the_sdram => zs_cs_n_from_the_sdram,
      zs_dq_to_and_from_the_sdram => zs_dq_to_and_from_the_sdram,
      zs_dqm_from_the_sdram => zs_dqm_from_the_sdram,
      zs_ras_n_from_the_sdram => zs_ras_n_from_the_sdram,
      zs_we_n_from_the_sdram => zs_we_n_from_the_sdram,
      ENET_INT_to_the_dm9000a_inst => ENET_INT_to_the_dm9000a_inst,
      clk_0 => clk_0,
      in_port_to_the_switch => in_port_to_the_switch,
      reset_n => reset_n,
      rxd_to_the_uart_0 => rxd_to_the_uart_0,
      rxd_to_the_uart_1 => rxd_to_the_uart_1
    );


