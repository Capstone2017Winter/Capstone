��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނ��>�(Ŗ�6�eQ�d*e��!i�v�4G[�\)C��S� y3�Xv��XcϷ�z���B�}��uE�Oz��q��̷s��n~܌W2����C�x��.ם:��˂S	�J�����ڐ�
�^ �	s�'�%���gM7�� �7���8�߻�So����@��>#�wiE�]�Da\E�ʙψ"�՘~z�X��)�f��D�y&�-��8R}qI���=-@Z.�������&�B�p4Z��q��M��c���j�R���AFW��\�T�Ɏbof�#<Y�^��c�=�|Xi�/7��� �#F�	Z�om�&��0�^�Sி��hf9�.����ѫ�v$v�������'i�{�١��! (����B��@������sl���[�df��sp�R2���*�� DƝk�L)��,*E���Y�r�5�X��9��d܈Ʊ�t=�����Á��ݺ*�?�1[A�c<P�'�c�<K0':�R��vu���l�q�'6-���a�{�cG��GF���т��Ю��s�"�e��b>ʡ�c�#���w��ϗ�W�F�\'\��6�#�2O�ghnO�]�Q[��v0�	���P�x�H�N���j.��l��O[���>"_.�L���0X���,�����-�帪w����;�.Eϧ�m(�ʝ���{��0��v ��'*Ԫh�(`���@�E��W�||�}�������*)�2�˴i�pF*e�W�TL�H�4��ۧ��kJ��щz�\�p�ࣈ��q��m�R�ϳU�K���k1k�C�c�2��ώ&��M�ԉR �h8Nʿ׮%hG���MTm�(ޏ�|���44�wC�u1�d� �&���Ì>j�k��:����H���@������K��ˀ{(�o�*
 �|��=�M����WF8b� ��M��Ⱥ\�T��^�|8�&�/�'��G�i�D�e��N��e'�-1��˞� Y��7V�)��v��ǴO��ڣ&���U�\�Y��ƿ��O�r�y����OP�?�Z�u�p6���\>/'T$���i�[���X�gH���[�р� �������^��$�	���B*X��̓�L���b��+�ɟD��}�l4V�qOB��i��\�Ѣv�|*��ٮT��@��+k,t!T�[�]Z���Y��{Q�G�r��0�����(�.��Fq�8�ĕ�X�+���vm�����-�V�u�>ݞ�)R���9CmF�5�>�ug�#$���p
l�m�>���{�2d>O':���<��{捯����Y(�����d�d�m��:�������I��]73i�X���d�����D?��+�(4=���j+�GT��P7y���QG�y���7�S����}�5Ed!GS+�x��}�Z����e8c�rk�c���8�D'�!�Է�)�SX:�7�[��с�P	Wo�p��80�˫�ȩ�S{bO,����H	���Hw^+��扝��hB��;�j�}sY ��c���^�Gn0-����s��b��c�\?a�%���o[���p��c��̶�{����Yr�aY�GE�&9���WZ�����l���'��+��_��]���ż��$�٤^�����F�	��i�Q��|L(3~���]�'6�P_�*ɔ �)�h�ޮ�%�V^��L��c�p�^D�7�':<̠Q^ߢ.��ң8��K�4T��ڧ71�f��CC�k\#y��ڦ�K��<��ng�����Jw���tG�S��C�a������5K�V+��z��l����Qx��ɵ�㱩��
(L�=��T�l\�f>	hu����h���-�]6��w�{�!�c��h�)���y�����~A�ԯ{�ޏa�~��)�����G�h�p��0��@>�w���$/��~fGގ�O'�X�"�Y����������Ի�BW�g�'�,���A�̧SX��Z�l��u�����^`��mdyO�#�+�\u�ߎg.�P,�r��&V��h�����-S�.U�8v��|��\�U���_KB�����j�)��冄���d�_��)�����~D�����s�s�_�X_�.�h8���!D�r�(�۪rY���
��Iv��"����~�5��!���|��h���P���L٪�\7�X��1��s�1d4+����h�@mIh�QmF��ų-�8Y�[}��S�Q<Դ7G4�W ���*�wu�Da`��qK�>�	=�d��D� t���
����E���
�?��{�%S��Տ?�tz�[�;k���-!��Y�_��Z85g}��9��R�|ذ�����vw����Ͳ�u?>�<��l�������l?�}����m14&�`��/����r`�t?���G=�p%V_��I��y��Qǀ;�4�6h
���c5��S�lq����<�����jt�E+��{���˝�C��i�?�S3�eϲ�C�U��R��(��`l�_@�I�ZUn��R`<��o\E�h�OO�qE�"$���67��*������"���g�ؽ��S��������P�7*�?�8l���j�)Ps@07�M�<�<��dB8�a���h݆�h��R�o�V�>�S�OT�![/�1��~�p�oMi i`���Jo�"���@����oc���ʮ��"7�����J�F�w�ð��<�U�C�cƔ���|o�l�H�7��d��]��I��)����)�3?���FlJ�o�����<�~x���S��Rh�g��L &�A<�Mʆ��F�y�����Z�L}C���\V��ɹ��2 �⏇v�Cw���xH�B�=(����Pl��MQ!�d�|��Mec�gDz@*�[���ƣ����}���gԓ��z1~(��mJ��k~p�cf���]�W���)�V���ѻ6�lk����u>:��,�;j5�ÀdGÒg�:��r�I���JZ��/���E��s���\��Ί�������.�0�s�t�YL���+ΈQLtE�kc�g���!0S�M�H�L� �����r���]��6ު"�2<,�`�����W��!��"���]���]
=wyl\�c�|�Y��h��~���F.���r�$'�_��Y[�(����������J�yI,h%�h(�O�?�Zm4"�;O����x����u��>��S�c�ԟ\�;ij:�"8��FWȦq3��U��*?�D���j�3���w$�;GF�~fo��`^W� n)�8L�;>Ŀq̠RxH���������������h���K���Ҋ8�=�����.hI�v��?y<���U�Z�|' /;�$Ň:�7��/ ��%9[�0ˣ�rlR{�\=�+(>��Q�^8�DTg��e��]��ʸӝJZg��Lݿ�A�ʊ�_
����MՎt�d���fPb���<^�(���߷w�9�+�շ�]���`T���0S��I�y�ݶ����_^C�;�'�1'`6�{����)��ρ��F�٤7��hV�X���Qˬ�HIɘ2��W���Ҟ!&F�	Gl��g��ƺ���"_��<�Py�8�)X�I�	zD,a�%I;����|�����M����)._�l�ձo��������*���	�w<�{�O:�G �޼�ظ��Ñ�3ֳ��mڊ|����Q06��"�xo��h�4 ���6�2�m��2�"�PX����ib�����.�Cl6�Y�T�E]�ن�9ɋdD��^r���5����$���t���0���2;�/�c{�b&IS���Q$�М�O�@�uF @����V�U������Mb�Cj\xw���*o�c����tN*�œ�������Lp�.�6g��i��e#�ҲDt4 F����>�娣�E��kq�7b�f�g�J������C��8T)lU0(-�@�E��:��������`�;�1/��]��j�Ҁ�R��Y�K�zA��ݬ%�L7bTi�%�h2&�����jƩz���x*�����};����=[-���L�9�Ϣ��V!��+`9�g^J�v�%�:]�%'�Ip
�Љ��k�V��$'�57Yq:�:���c�k���%�c��6�Ypl�� GFe��O���*��M赌f�F�W����U�>c�Fh�I����y���%�V\��VA����A�4���D0���N��,`�ƛ�����u��������1En�>i�T�s�d�N���v4G?�(�d������]���B*�Z��~���]�J�V[�����nO0���Tq���"�|���F4��\?b�B+��U�1�LW>���y�����<mvHK��Nu��=e�ˢǦ��
�d�	��K��}�D�XGEu����
�,�*k���S�~�T���z�Prի`�Mљ}�Q�̛��k�戺R`�����}�[Cb�W��{X˽��Y5�xP��KlU7~8|�L��<��.PW"/�{g�!E�1
�9I�1H<��/J߂�l���'�!8���NVQ�i�k�Pm�3L�`����:�,�����C.8�S�����E��J��<%Z��%�#0s#ۛ��|�L�$�M���A�Vy~i��`Gcg�<�b�	���dzU�ӝ뎣�+�:Ƶc-�ߡ��m���M?C��s�7�����E���2\��rF��χԸ�*�?�J <r���6�ٻ��bw���H2,'��wF ������m���aߨK�������{%lVt�jA�(����&T���<�]I�6�/ꄒX�}�i���#$�!lBj+��ڑ?rr@2�������8<��8t�BSj�i_�������-��4�+:���`��O�lt�o���{n@RD$�?���~b��:ni!~Q@͈vB��^u��;TL��S�5���	�Ng?� *t��4�Zq��2����h4 �7�{L�9MI	���_������+-b0�L#�:y�c���ojq���6��P����{���L���-k�	���*��C�Ӽl��P���G�VBqZ-�.	ᶕ��%����E��,S����<��.��E-�����?��Śjvv6��iL���i�[t��Z�178�����<�%�4 �F4��걡d�>�fqɒ��R��x�h~#�X��?"�=aV5���vm&LJ�K�gh����&Z�1xh�f�f0*���1�"�.`#��Xe/]�,86�N}�n1ј��sf���O�P�7#,�D3G�:!A����|�[����!��	f�����@��ʻ����ؗX`~��l'\�sB(�eG<�opȄ���v_��%`Z�>e�G�ŒOo�t�S!t\�	=-2������{�y������uSJ����e�s�#K��~�)5�"�$����C��|2�9~Qd����icK��Q�r��F���L���K^MVEWLR���G˸e顣$�$Z����ժ��p!�l��;�	b���;��ԟ$���Ԝ����R�ެ�+ߝ�l\6
ǃ0?֣P���{���EY������X�F�@3�L��b/��J�^�7���h���@�轅���哉Z�:��% �ہ���S:|gîD�K+�
���-��vr���w��*ק`�@���(U��m<����D�4Ɍ�>? x�
]g7�Q�)�}�)���D�r;��
ȍ�//?�>1/�& ��KR@��q"�٢����N�{Ϳ���!ET�����;�7<bȫ_.�?WE����E�l��B���Q9�p���E᫖X�$:�=R���1������/�gm n�XC���"XLV��^���;JG��D� W��GW�{��R��K�R��Ƞ����XbR;y3�c��NY� Dj����[���Ҟ*4?����G�7�0�B���P���{�*s��]���L�5�p)|�B���d������'��qԑ��	~�ԭ�k��U"�)x�3�
t�A��d���qi ����tb��{�����(G��r�����;V�Z �OJ|(-�KEO"�m ��N�-;"�*^�ՀG��w����ĝ�����tm+�P��������	�X=�^��$`�M�FS��\@+3-�+(v�zn$���w�Cv�_���H�������˥�슅�����yw�ﳈI��^���ѕyw�l΋�s:`=C�
~�A���~��>^�"�6%3O�� �������1CPuK�l����3E1;`�@��+�}!]�W��|��,�!*}�K ���o�'���_=k�"$��q�$nO��N|��K�7��jΌ�zDRW^�TA� �h������,p�4!�'Y����}9/�o\h�v�7��x��b�e�j�<.T���$�I���\Q3���C��@4&���~���B�g��{]ۖV�D�:��g�c�/���&Fş|���� ����e`��o�L&b�k�ӆ��ǽ�sdHc'	��\HDL�}� ~GI�(
�$6��f5+�}�+����(�bXJUp;F4���)H��
��E��ľ~y>�սz���XT1�4�X6 C�k���Y,t[?�p}��0g6|�����w�X���a�7�3ab��&Ot�Nq_3:��R���k�*�,_��51�J�m<(�����
[�M2m '.�Up�)	_��fE}|�p��O�I�ʨG��J�x6A�\!��Z{'-��eF��q��>k�f�媝Ad��u�>��A��(F�
$��;�[�ʟ��-�4;��&��Ӻl���J7�Q�$(��B�
����F=X'帗�n�J�Z@����"�'/��z�����Қ*a�E0�-Mp��rfX=y�/ȋ��)peT���K��2�n�1ЕF/�x����u����P�UӼ#yJfΜİ�� �eMl�P��=��5R��XF_ 0�\��u�;�8�/�)+�lt6p\u�}ҏ\����P��Z�t�e� 'V����Ѐ�OPW�--턉x(E����j�6Nve�9�����Z�(P�`�~~�p,i�C� K��[)�m".w�ɺ�dp&jA�A˱���;�W:Ϣ�����`�!�`�Ѓg��?���kCųs�0�U���5IHg��8'c@��u��
�V��鎔{�<D���uE�f����ѻ�1�Ё'�3�wr�,��d�a����C��G�ݗb1�G�q:FB��y�0
`A�����h��_n�i6�	��e�߯"X�%�W���%�5�6�hm�N^�}�$I�A�b�����k�p�n��"�'Z�XV����~����B``������lZ(�NK����Vԣ���/Qm�j<��F�h���Ǌ�����`ߤB,z��FFF���T�,� x7"�@�UR��&w��Yd1�fhf排����9Z���jo/O��=dݶ�Ђf�����	5;R�Ǩ�,{����3�;��5�a�ȓWu�rACm4+�����pR�� �4�ҥ"<��a�>�5�y<�brl�[x
Y[�y�&��a��������A��)��@�-U����7�$(I�k�S�yj�ϛNs�����'i�V)�(+Ƀ�ñ+���Q�+�+�-��s�2j��$�!����F�s�M�6'�x{�� �/H�z��%d�T�p+TF� �}P�Ϻ��A���l!�d��VCž��9�L󟤅�����o˨��Dwh� L�Q������C��)���j�lkG`��EB0�'�|�=��=�*4L� ٩7��մ�j�^u�`�(�@Pʃ
�&�Sk�� `NΖӡ5A�;s[oND�6�6�vN�;k�=)�.ڒ��p �� ���zZ��u�0S�KGG��7�ugY����f�c�1¶�>�q����Q���m�\J�����UE���`�2씼U�v�]����݈q�h$z�3u
�[���D���� ز���<.9fr�}(�K1�}ߙ���і�����'��-�ڽ|�U�:�EVl�*�-�إT<�΋!�>!�����R��{'��N�;<�m�ްQ#	�v�r}@�	�6[�u�	 �Y�s��O�&J�����M=ߧ�(㚦�NYff��B��[��"�F(!��j�����z�	��&���[�}L鼢�jzb���K���3�|⑔�1�Ӆ-H��|�T�=ՕG_ӕ�R�m7��<*��-Sb擪�U��73ǎ�����&�q��Ŀ)}�$����w����,F^`��kK�h�� 9��
�as�J��	?�)�o�jXr6j|yY�H���7C�aI����(�*R`�D)(�wLЅ2��ލZ�P�Vd��m`���#[x"��؋��0�z�uZ=&狅Yb��RӚf;�_j'P��B���0�e�C�L?j�;�]t��������=M��y�t�����I�f���ڱ��0�.ζ���#(����/3��)~�� C8��q���̃��s{F�J���ӱ�n��6է�p�#C�XjU1y�oo��
f���h���a�P6�H �z��)p\�v"�K��	��2����4��b;��]x���F���Ҋ�z�1]��j�`�]�rG}�)�"7�?��B�����l\#��N ۘ"1,�����͉������}t�/�h���q���[L����g)�)��V���H>8Q�l�A�q�Z��j��+R>�Z9:�x�w/h�m��'DT��z<)x���Q�PS¢'�����/"14�7�`;���^Ŗ���!����G����Ul�!1�c�\P9b��L�����f��~�+�އ��_QQ�{!�ԥm�M�'=�s��C�)����k���d���]�5��ymE�_vDi��x��o�r˗:U�sq��w����v��Mt&�w��1s�
`��'�����|���?|-QD3Ɯ_R;�FJ�1�l�$��˙}���\�N��l��O,#@�����5zVۣ�)5
=s��56V�&�~�P��ƎA��[�d�!�Ӥ+(�S6{��
���:B3�9�{���?"�?���}4sj��c���(������*^`W�$���.������<�p�2j����ڤ�4���aĬ5�e.�0�L�n���m]d���'׊lǲ��C�s�����p�kg��伶�U;r	�K��&���օ�*I7��5�ݓ�dGʈ=s�( /�	%iZ�s�>��1�f�H�it�4���<r�C����ṂRP�T:͝�����0üo�0I#_���)I�&�e�XSy��s��<�
�E��V:���O��d�8�Յ����5 /=�PE�e�9�uHZ*��ȭ�_��E�@h�J�c�/w��0�kMH�̙ky9xvK�ic�nl�~�-s@�E�#�����;g��0
�	j�x�Q4ZM�?@�6Zx��@=6*�߹pŅ���|As/~GM�=9��nW��X�UP�Է$w�|ŷߢչ�����%��š�2FO��~<~2��	�(^9�ּ!s����ܠ<IDjX($�V�`�W�>k�%J8��&O� �M��|�S�Sa_3����뚇7����h�<�Ȇ�*_���F�3�>'��]_�o����-\���b���B�����⏷t��El��3[nC;t��̓�"Y�;�W������Pv���/'�`!���#qz�c�Ŗe_?�����ak-H��	f.&�۹��́���=� o�g�Ϣl��ܬ�rN�����Lhz��pմ��t��]������ �]�\�33�ه����^�Z�>������Y��|;��lMT�#�&�����t��X�9 �����kNn̍����*�m/^q�)=GG�\�,^qdG�\�b�����4�fp�	1_�%/��[�D+���ﶾxD�((=��,&cd#�n˕\С�n	�W���{��m�������zMW�b$�k��2w��,�M��{��Y�ܵY��"�[(!�4>j�W���iȧGv5t��I��%��*��/UY<������jg4ח�j ���?��������.a&>u��dT��f��ԀxnG����q�i�ݸkx޴?���j�����(��N>[C�t��|�ű��݃�0��I����+wek*�[ǫtHLx�W�eͥ��������:�S$���;�N�_C��r,8���RP�yS�%g��"_��&t�ct�f����`=��_`�ј6�v��W�z��5;���~J.����]$�!U]����Or�!���)xc[%��Z�H3Z�"�DJ�D���\.��ܩ1�`���e!�|�*#x2��L�ho����]$����ER����":���ߢcY��G����@З>���U����i�A��r�,j��!q�i�C���z�wE�t N�g�!�zO"�"����T}E[���e�����/HQ�#qB�y��H�:�*iNx֔C�`�6��>�B^�WI^�fV�ٱ�M�������+;b6���ȅJ�Uʞ�/L�g��A�w-�)giԑ,z5Z�1t�#�s�2>��[<NE�c��?������K��`<*1���o�L�k������=a$>1S�$����%CYf�y�B�X9�niR0ؓ8�
�3@St�;C3��@3���/�E�ב`����lt�&jb��h1z��/�c99�d����Y�u?^Ђ�O�k�s�q{��4L�����D�����gtm�� ����smY��3/း[�&8fL�%`��+"�[׀^v�g2�`^AX_�M`�C��;Оѝ$��s9tw�Ҩ�q�oc�9�Qg@�?W"2��4�'��;V������dh��o�Mw�;~��n)�"��J���>#i�O����Xݫ��"�DW`�Ղ6�T�rf(�_��L	�R����I2ψׁ� �h�O����g=���ș\�#�} �L�n�
�hA�7AEQ�����6C/!�F/!p��	r���FEL���}n�a|�\@PU>��~���x�dg��
��	^h�y��*��.�����/�ҫ@����C��Pᢃ�/�.d|-:b���ނ�eVt���@I8��� ��gqXb{2�Pp�묈u-S���9��#*/�������%�!�+���O�m�U:�`v�2R	(&���L��)J��-ڙw��=b�q�n�ҽ�n�X��h�5�ܰ����L0x�k��c�rA&ç �7�[#$(��(ڲ9u���&�a�;�Υi��?U�d�3�p��P���!�g n�x�1F/��S��3\��j`�.	Tah�eO��Ud�"(x��Iͮ���+�R
.*��	k�K,5k8ɧ��߬������bI9w�sW��u3��}Ľ=��>y��M�_��b6z8�}�	��z��v#��@��% ��;&��������Y���Ki��s  '�@���.���9�BX��oV4~�
|#E� �z�)��5�k=����qG��5�����n�1��/)��G�"���[�H��@�s�HzO�듢@�rZ^Oq�$܃u��)9�@d�&K�u|c*w� �	�C5p��JmM�r�z�Z.2b1���t��p��]lV<���K���V� ��@�d���pmɉ���ը�\x��諨�phk9I2�(58e���i_)[?2-N�8.0��W6�T�T�&�Y�IPD)�򠟧7�D�EWrT��@H|Kte+h+ĠBX#I���.����a*R�GӖ*MhӤn�N�q�U��VѾ�:i����#��ף�7�6Z��o�<�ؑ�]�
8�v���y�b�T��������?�\����[�����2�kVe�8�̈���?�ճ퉻�5�h�_�γ6$�{�	�=b�`��Ƒ���t�hѳU�"��X�Q�m�bͩt
iw���|�����ꯩz?��x=W1�)��7��%���?��}�%�!�[��?�k!���7�`�Q�ۖ�]������C�����ر��K�B?Xx�\B�A�nu;��,�"�N`9UH��gu�kZ7
��\��$d�l��s[��&�qݩ�8��Wx��#����H"{Pa[��v<4�I�Mǰ_D�
��/)9��mF8:�3�H�'��h�����J�]E� �V�N�jP5:yE��3�9����^�#B�y�&�Ÿ/���>jFv���NP�5Oڰ@��^�h�B�`�a���)��=؇��B���񵷂�E��\t%��k'��l�O^)ׅ��V��Q��w��Ao�aO6#h6YR�5(����{���N�\w�>;�x���ۣ�Z���j^��Ć�	LAv�'9�ʋ9��;�|[ܻ�Y�@�8LU��yވ�8�]����6��1�:^����\�d1�3z��`>�S��0C��R�P
vv��'e}XEPmՔ+�r�1i,��Ǥ�H�i���@��TUb�ޭ����WG���w?��MG��KF
�])_Sa��T/p�WI�3���r��9�P:��3G���;C�Q`��������V���"e��t�iv�jK�Ve�l��&
pfC�n8�ǒ(o���D%AD'5����%(M�㌳�ul�G󙶃4�M$%�5�����9=�3��;��\p� G�f3�G��������7���ӟiL �i\���k>~������OR�0����Y0��+lִ�a�<^�Y�c�+s g����'���RG ��!�~k@��|�~�d	�������.�����c�/�h��O�/�7�8BHR3�N�K������;�Z�s>8��w ��5�=:�Y�{i�v�uCi���@}j�j�����h�$�}������L)�$]�;���ډ�8�W���˼��V�:>�˙�E�А}��U7=FN�447�b��e�1�ᦡ�u
h��Z�Y���_���Rh��va�}Z׆�x�C���51� 
�CZ�]�d;�W'w��2]��6{�%J,�NǊ��x����?�ӂ?�}#�����6#kۥ��yD�r�[� ����U����o�׌�_��w�]ť��_1�%<v�r/��R�f�n"<@�QftL\��I�;���2��Ũ�f���~R+~���.�g
���baU�<�&v��)���y6�}��X]�P�U)4z�OrQVK&�0}�q���O�����q]	z�cʣ@�v�%�L�D��"�ޯ|̵���?��G��=F�%���n�������Tm�h<(Yw���/Ҍd5|���_|���F����S-����!IPg�^�Us��8�l�5�FK�_j#8�#ϯZ$y�%�ǣ��5zɍ�k�H))�G�W�jp2��ո�(2�=�3�m+7^��r��3~~T�FD6��a3$(�q�)��Z�f������Pʘ��U;�u���6��=���ޡ�\�w�'�ٟ�w��z�@��ۛ"?z�mqZ�P�ny"x�
�u��/�� 6_��'��ox籚x��V�S��8����Nr؍�!��! r1���%�؉ݵ��V>�^�����7�OS7��Z��@��ؐ��E�@�:|?���W�15���_V�p؉������[��0���t���6C��%n�
I�����*���=�c*O��jI T�G����rͿ��J�jY��WU�)��"Ӵ��BԦ�g�6a���X�ّ��z�^��T:�������ȇ���o⋂�Pu���̂r��/M f����X��f�JY�BiG��<�(JYv4��)
�����BpA�-lI:�ְl��%�W�rIe���5��d�1�)���YH	AM�PK�щc�.�1�l�@8=���E>V���)���L���9�̅�h��|�]�R�-�z�{Nh���hA��Mן�-���4����mƂpP�hȩ��#�iU>I��y����@6�+C��a.��5'B��F�T<��c�q/E�1"; �ې���s��d��/U�M>�m�N��M��� �w��طW�<�X���}��~�;�����*��pQ�n���S���G��G#n��OC�� ۬�?ь��!�{�f���qo��O�ꚋ2�a�J$�R"���t�o�<��'���G�t�ˈ�Lه�}�׈m^��<qk���f��66�xm����pL�m����ː�.�֊y�;�s��"��}��7&�|Be�+Y��Q�DEA��n�!D������pY+��K�z�W9�ɑZ䧌kK��SkFDO'W�y�U
wB����uo��kXo�=_��tɒ.�����i�=�+_�����o�e���;<�*�*8��Q�	�&��S�E4L1(V�X	��ԅ'0��VeW]Q���/�؋�ݛ[�S���|Ak*��$��ź���-�6������RV��NuJ�Xqe���Ni�c٢� {��n�@�i��gRQ�#�F�T��@�=Q�._�i������'Hb�H�)&�N���z�0���T�EC99��V���.<��M�O�{��@q5�a�'8d��u�(k�5�c��5�Ŷ�@4���� @Ū�����q+�5�v��iT�&2d
��c'/����9�!�*&���$�1}|��Ά>Ǡ���~�V��;qc�9h�'�<G�A��$7� (*�K``��.X,K��V�s=7�9v.�`t���T.=j'��/k~�����{�8Y)ŷ��E��;h9��w���1ҹIE[���v��^q����C}nh��`��D�~]�MP���/���c�����Y5��"X
g��.�ݱp����{"�����̣�{l_�¶�����`��.~1PN¸��G�Ryڕ��"��}�PH�d{� �S7h�Q-W�tj�"C���	�G�WA�C�R a���}�2LڡI�5�;��7�I���2 �۷�X�І�N��%!����0�}�`µ�Y�������S8ԯ[�u�:W���,+>�ņ4N���^.W�V'��t7�u���7���A,�?V����n'�%Ы�N��H��*�؄meh��1PP"o�d9�E9���L? ����kz�JT�	���&2�}OE�V6�wK�&�.�5��1���{����}�
}v���5��0"@_4#m�!����u놮����2-HVn�����Rc�J.�#���6��G@��|'|uarX�~i�c��Fbŷp���fK���3XdQjb�#�
�M
}�����
�� E��?!र��1+��	�c��F��`�{aZ�Dd#���TV	'�2��$��L��P��u�	Aoqqf����4,��g���9��f����y~h� (岌�g��Y{}���noc�1�t������f�-��ܿӠiW��`d-TV����� B��r�e�>�j"*�M�M;Լ'E1TIЌnkF����@Uh"ɴ�șs��%.�f��0���X�~'�ON̰�`�4��!�­�D�2���;����)����p��e�*b/F�d��F�{�����jsQ޽�Zq����keV�C�n�-���O�tE�FժK�>�TYb��i�u�`��#�
Vn �7rB�:j��D������nY�{c��@}�ǥ�_sٛ(�/3w@'F��63yc#K*�2�5��iA~�'E��H����B/�;!��$�EG_����F7FR��xu����W�����e?H' �MѕB�����ĥ>'�N�	/G��16�7��:�ʱ�����Tx�r��-g�?dҮ��Y��:�y�,-�ל�ZX���۲�&�]���������Y���ؔd��hٳ��w�P���fp��A8،6y�L�r�����[�}�n�<4��O��r>S톕a�>.�%m=|�E/�+��!(�ܪ�zSe3[��Ӕ;��P�s
��gjȹ��nq�h;��UY'��]fsl��g�����@U�4�IK���V�'rס���@M*�! n�?Ƥ}���N?��^�^kj-��3�!�E+��E�3��Kc�?l�=}U����{ss��S�p��٪�g�o��g Є�}[��� n����3� v���H��B9%`�$-ՁP� P��o�̴��/��o�3:�Z�ЁdA�rlB�Y���@��}���2�1,`��N�&�jAX�ԣ޵`�`�h��b`�����%2K���t%��©�A�z�UI8:��gru��A빒��7UV�j�V�s���]=;�����5a|~�`a�^�����<i�b�?�8��hc���i��ӡ�KI��d0U��������t-�N�Hu�X�͝����a��j9�JkOZ��h#m�fSE\KJ�e�mɖI�u��b�����0dl�7x/��о�^��CC��m��
N��i~���a��-k��85��j�
�N;\��GM5��w��M�Q{�eW"��l�O(^��=�{�_�����Ά=��0���[����7!�C���7D�o�V����\�U��>	b����xD#"B}F��9�TЈ�Ȩ�Uz�^egY*`3����l@H�M�L�����(�lʭ�I�S��f�/�V$����8]�&R��4M�f�[y?�X|�E�H�дN��:������n�=��t�� ��~�1���sp��[坓>�cp�c�_YET���X���^�@�(�l�_<�:s"j��µ!C�~�e-}�A��05����'���MG�DNZ
��yr$\n������{l��ph�Tr��A�,P��DJ$�%�ug��@�ў����BpW����0jy\w�$�,3�QKI@�|�1F�f���<0d�� 	�q�6�5�+��9�敻ս߽c�
o_�
���I}��@w��]I��W�x~�X�c1�ĩC��[��0����_x-��w����*�g�6H�#�(8�<��o��S�,��ӌ��}��ao�>T$�!�I��V��JD!�09�a�[��.+��پd��/�o&�Hݸ:� �2�c��Qw^6��)kH��3�r��Zʮ��Ā�p�B5�kML�\���'�h:��4\�,p6�[�-�ݗD�aƿu41/���|L���r}=�x[�s����0Ly��5��8A��(<����+�v�"�Q7���-�0��/�d�R+���k��wO��..@�g��B�$�vm�>6��R'f�?��GƯY��:j1f��WG�HXi�3��Kۍ�*	���<������ڊh'�켲C~��5��a���x�2gqŀ&�"��ްT!�T��B���٥)���/��ilUa� 3#���w;#T�U�d=j1�o(�4��(����v=옅ڮ�n��T���ڱ�,T�||��KyCh�����K�U)(l�����Y�6Ն��&ϑ����}�K5��c`f�a��R�MS��ݙ���G�Ny�4�Ģ���Z��u_}��6����;��\���D9Y䶔����CP=�e;�$Ʌ��H�W��$�ە��p젬
��|^�A2�s;w�u;<,K����(0g*�D93R^	<kP�	Ar�4�]'��H��.��^~N��ACt_�!������%1��/7�HX�Q܃(�'��@�����$�i$�k�F���ɢ7a�7�M���o��\w#�ۖSV�%,(���oB�m���Q�hD'wNz��G��F�l�A�u��ӎ�>�!���0���C�M����	�`�����b���-��u�ijU�K�ù�
��2+ �}ҟp���SA�2��w���[yt�<<bZ��_`�y(�y�ES_Òly:(��Ix����g �r|]K3�����}���P�RD���3K�pn�J�I��kͪ�j�K�*�Eö���������	�48Iz��w|���� N��*�l�f���d <�(��db���xE�/��9ߔ�nI���������3��M����j��1�u�Lq�$u�`W�H�v��f�6��ޱd����1���G�� e�F�����!�"�!@�K�j�`��`���ҭ��cȩ&YK�}���⟘�u���$m\N=T:��:����k���y�R���3Nx��]�u��¬\Go���m�ّ\ń0Z���2[D�/��%E1/ȯf�(\ ��#g@�
���[c���S*��n�09�^ֈlͦ�D�^��oˮ{&�	�f%�SƘ����*��A"t�����ZO�/C��p�WVQ��"+�Y��.erQ�4�)|
�B��Ӓ��C�xl�b ���{֢��ii���?�׉����?��}����f(4ʦ��dT�gu�{���Ψ3Ҏ,wȌd��E$7���&2��V��t�
w��4��a'n~�N-��.��s迄���������y85��6�[�0���u��4�D+i�O|R�4��Ch�J��ʢ[�����Y�K(�O��+���u�?��Y�^'9ڀ��)�Q�dJQ%�8�C�b��җ�Hˑ�c�l�ǒ�I#�7:�3K.7{1�ײ�#��x1�X���*�u�#�m��萙�ߕ�ܣ���3��X/��w4w�^�l�+�3��3HYן��]�����#Vm�윺�֏_��dj2�a%�������4�ϢS����������zZ"�f5< (fS �R�9�pq�(f�٣V86R�gI0 &btG�l�M�znؓ��sE� ��˭c���s�-]K��M���g(C��5�\@�v$�����v�P�	@ߤ-%�,�E�d�v��^�~�B�����|��&z�_D*���Lp[�?uXP= @��r�V&BvNV��8}Fs.�oZ�O��1��q&n?�����	�!عG ��0�j���]Č���ڶ�mL�e�T�X�#�i����x|5��A66x12wFk����G���D|t�n�j-K�taiH!G�=����Cⅷ���u��8e:KZ���(I	/س�g�x����5�U� �Y�w����p� ������B#�� �u����tti�ŉ�gDT&[�6 �~���|�gd?�IZg���AS��V�WX��D�0o*i�E�
��i�����I����dw?�<��6�c9�!�ہ�Sԃ��� N` �"����g������J�x3�0���Y�D�HtZ��~�	5d��Q��[����X��S��:4IgI�E)��ͱ����۬a+G�o3��'AX�p)�9��tu��TH��*�ل��F��E��K�G\ub��E]�U�{�8-|1�C98��a�#�3-���ߤ&��mP��%^p����N7��$��3�^j�#�*�I)�9ޢ�߫��E����@_�Xw�����;w@�{9�/|`oO����<G;�c��񀵉m#�1G�+d�_���'�/L�d�����n�	�٤8�)�7 ��P�s��i���R��Q���ե|�XE$�xa�݃�����菿
[#X%Ǡ�'����f&4 p!�u�.�v�|�J���_cwI���o�D��e����o"uZ��7�
�������M���jP0�^S�zb!�cײ<ġ��6C2'[��c1<V^T�e�*�M3P䫱�@eP���"�R���J�́�Cx����!�{l���K�@�L�gmp���F�-�j�i�V����ru�?��~�\�ü�5JX>zL
���)�\����(3���n8�r���wg�8*�YRVM$u	l����?�sk"�J�_����?������")��5ߊL�&��i�+s��ͩa$V{a�M���Y��*;�qE��1�g�8���Pe�:�yAt�v��t�w+s �����
�Ӏ�'��=y2��}:���n�~x4����4�� -r��^��k`��U�B�%��Q�
��c�x��N� O����ꤶ�k//Hv�nuY��`x�$[~�����vm�]ԅ��U�û4hį=֕>Q�9�l)���J��'
xEhh9�ЫgR��oI^Li���}�3\g���+�E{�p��H��R��]��)�P>]!p,��5���V�?���n*JY����QJ�~mW�Cr��=ʹ�F�,f��D�R�Y�N��U���^����בe�����FF�&�0M���+J/�Ow��G����ԇ��C��*��\X&��s5�؜����ts4�_%u��v
�^C�C���b$? �>��9(pe�S�x��ő��o'$�;��u
>����������� �F������0�1�����U��U����]zgg1<��s���?���"��ڨ<�䡀�at]k-���$��gN�>���9t�N�O��rR���aHv2I�\.�|���eRS�W!����[�Q��#xUj��֏��ܤ?|�o!I�l����|�f��A2	u���#�fZ���sT�/�IO�kOWg��21���3˞���#L>��e=��j��aa(�S��I�ӔGǳ-R����0d���f�Xj�"A��E�@�Ց�6y��ڗ=�jD6�$8H�4F>�TR�Z�C��������{M�^z�H#u��>l��ۀ�Q�S�~.$8��K$�[��]N��ܖ9���7qs� �� ��,>��;~����y��0�Ӧv"��.�:���:!E�Ib��"w@��[�yĻ��Q�a�by��6��"ɠ�3��R��;!M�댏��o���A{�)�/��%��w�kސ�p3�Y�F�%����qn��
���:?�"�+
�����17�r71�F_����:xq�i�lhR���n�-��C�D~�XZA":����)�g��_>ea^JS^������ɶ�ؕ�w�^�B1�47�ZQks���&�����o�~�r%��YΆـ����#�b/[!��⥉����q�R\����V��"�¾�s�H�W*ә�$���E���9���^��� F���[8��©�4���W�Jh����B�[�v���@�o���T���N�b$�$��>Z�-2�?y7� 1��#�k��;��[�G��4��]t��w!�s��p�2�5�/Z�R���{i�$Y^����%\0e"qqF��W>��",`��s��
Ӻ�kqux?� �ԣ+`����n� I��β���R�4�"Jc�tv�0��*:^oc;Kߕ�RY.�5��b��n'���W�]����B�G�1<�*���j;��)nV��㇉�,�}��N�E͋^���{�w�W�;N˭j�g�a���O�Y��B�Ts�o���ν��ɂ���)�H���!�>�{'ݵFR��G��1b���F�h�X�
F�W"�$vt��W��DJ)�����7�]��+<˼�����ٍhe a��m�^Vdc	�[���TgV$�2�p�!I�n�DC�����ݻ�1]������sH&���y��n�2$l~�$��"X�,�?v��u1*N<��DQ�����M�(��vQx�d�W3u�X�x��%I�%�(����qC,zʡH�K�}P`� V�%M��D$�(*�z�E�eq�=%K�O�.�
G�)z��j�h`]�zTA���;ݰ@�9��;��u�{WRǈ�<�C4����!�{�u#����)�����΂��^� �b�Ⱦ�B/&��v~+4u���9���Q��@��Rqx	}�}a��uV�B�����	h�w��Z#��r{�O�f�u/C9��g�W�!u;�N�@+�����Jo�a��*���wY�����-�#!3}X��R­�����Щ�>�O�;>|���`%�����I��sTI>>8�xk����:|�(�tMV�?K���Z]�n&,Uv$^�������siu^e�i�jtF���B\�{^{�>�v���o��|GsW�(1�bLu��b�T��.�K�ěZ�g�hg�"�J�.��l���*�7��:�&|�4ڄx�5!�E%������F�[�c�]I�(
�^��q#�l��tnx�?�a�P�T���.�"����r�����h"{k@�����ء���#A�Y"����M��;���E��󭙟��Q;;﷗8��u
@Y�>āo�G08��s= R����yy� �Z������pK����6����F�����8��k����5�&� ���)��Ԉ��El�h&B)��_G�T�������$�#ȹh��.Y��U��T�L �H�NVT��Ğ*�6m�L37ɳ����H�d����E���{�п(P���ͨ�	k�B2y/=(���YBq��4�s�p���$�9 �
��&�7Mc�]���0��G��O��~�*���<]|��uyd5o���y��p��Ҁ�;姩��.����B�	��ds��A�L?(j�sJ�������_)yj�����b?:���ґH��T�8O�嫅j���ӴhM��I�6�>�劆̏,*�#�5��ޘ�7�--M���$��-��D���y�p/�؎lD�"�(��QlR��i���72~��Z�}7sY f���3.�~Gy.\r!��(�	����^A$���p��JĪݍ4�KuB|NW1Q����0�~�d��:�)�Y���);~�fD�����"$�!��5�`8�9����&9�
Ɨ�/�v(����St�d���Š��Q���NCr]Ì��e���}+$�����r�g��.Ud4����^u(���T�LA&ȴ�dA@�j��E�:��:W;�6oR�.S0��O�2'��)�2@j�n�p;���R��1�pDHpM���5�S��g$���lk�v��8\�_�0p \5]C|���	/��l��k�Y�mj'55]t���~r�=�=]�p�ј�˗���x��xgyFF.�4����>S�.��/���:m���!���*ȉ�L�z=Oe���(�!"	1�-����K���b��ό�=@�h��k�z��v�ZmQX�>�Eޅ�䓇�:R���i���>LC������<|���C��,�ڰ��fO6"y��y�ʉi���e��{<���1F�ǆ^3���5�c����]��#�Y{���@j����&�/�ä���F����kf��>U3�YZ׀��2=�$�Jw��i5Jbԋ��ȁ|�ۛ"3f(�I���.'��J.1ƀ-O����$��Xr����|�b���U5:�X�FVh��������z�=�ö́����T=�o��n唣�W_�U�y�ḫA��q�l�sk��}^5Y��0�#�uVZ�J�/�v;�A�c�����_�2D�(o�����g��������A����˭�F�����ww�]�2�)�j�C���+�[&�r��s�<&�doF�����J���D���iz�&�(��+`����F�7]f	�4�dC���*�R���� �7����_��\V3����`���\��V7�x�ŉP��f��)�}΁n|��R�>�c��'hU�Rv#�h�P�Ơ?|9U���Y�잳��D:_ضC��
�V�. �PN(,b&hM��å���җ��g�9t���a��3�L;؉٨�B�N|(��p>��͂��%$�,�m�8>�Nu�M��lB�w�~��}�Mg��d4Жףf���4uD�4�����1��
�â����˽#���C8B��I��R:{��pJ��M��ߨ5v04�C�I������^H��\�EO�(��#��.V��s�S�p�����]�H�N���!���u3���g�bC���<�Y��,v��JR=�m�W�)���Z�����N=Ru����'���W�0���)HaH2�\>`V�ԩ�үw�2�N,�V��("Oī��;^t�#z�Y��}!L)��H��GW��5���*�eL�E���j%�jI��f8��N�ܶ
;upPݗ���7��6����!�4�(�)���2mG�13R��&+�J�k&�����ָ4���f�'�O�	��~Ä��Wa}|��dr5w�R�k���G���TL�������xeG�
hO�2� ��9�8k�C�j`� ���)?e�L��KC��Q��4p�grj��	6R�
f��;A��6�̗Ѕ����/���PI�*|�"1N�Kt���k�&~�Oj��q]9��C�ބr,�h7�Z{��ʶݔ���a�̔����Y	�������� q�dɐ�H�V�e��[6������Hˊ�-0;��lk���]*�\�J���j_3w��/��l�#��4`�0Wʵ,��$�X�@�3�R;��ApH�w��O�Ś�.\W�z��4Dn ������m���h�s�,±]����-�Y��p�CX���X��IKevL��:_-��9��A���&ӄp���7�'NjM�rs���ݻ�$�vi2.�9��@����P�O�X��\H�fd���˔c���}�{�]*���]�l�T�+�1{x�u�o�6 R�\Ӡde�'-M����;����]\h�2��v� <ވ%�AP�G�ϩ�E3�o�?FB��������6�vj�Q�&��e����Y-�X�����a��>M`�E�u���P9�?@�����KyD�@/��ovqw����V�;�
X+�P
J�[�v�o+L���?2�À|����@�]�ם�ϙ�� �j����;�?� �R�$((��-�8��j�?�Yԓ�sB�]mU��&�b�o��V��H�z���W�o�q%���:��=�&y(���t���a�w��h�Hn;���='b��`O$"+Y?�d|��h ӥseѽCu��ޘO򳎜��u+S�d[��7ׄP�픅x��*f��v��#��X!⹠^�%{pQd/䢤����{�x¬�
e�D
 �g��[�e�	hqd�q6�k00�4n���i���?�k��盜�c�&���xε�q�Bm�8OGl�:enۨ1'V^�(���Y�פS-��{���&��Hz����fIU3b`�p��+�k�@�%[��P�O��Ai1��f\N=�����зʚ�
�l�s�Nl�.��RX#�VF��r�h�֤���CH��V�=T��ecv��Hg͂����tƹ[�u���j\p��r�?�}��[��T&Ǚ��BEr��� ���v�
�=��s��ͅ��W�_�%)���߻Ch�,{��TiE�ĸSӉ��0�RH���L���o�>����$�a @�|^E~����!
����4�X���@���,H�{ʛ���01�1;
�5eؐ/�Wӽ�Lh�>��7%���Ұ��
߳�h�Z���t��CB%�_IT��.� 1=,p.���*ˬ�=n,Y�w�*�L[x�!,�2�x3;Œպ��d��$@-z�NďhR$�MXv-�l�
��-E�e���E\OY��� �;�Z?`H���{J�e�[H�Nn��↏t�}hi�2?]�7�}��ՁP�Sʣ��q�7��13G��⇫�
���!�>��3���FҺ	��{��
:�#9m���+!��ۨj̨�6Tw}����6�65\.����c|��`�m�OU��.����������cI����}��r�G�hڹ)�+f�m\�}p���i������^��ny%>�����޺jHн(�4�h����91�G>%���9�~�;F�q,�!=����v��:�oe~���ir.�Z0�#<������S�Q�vw����B��ș[�Rp�|��V�����n��x²�I���q����Ʋ:R���0yhB>K��e�d��� ۛ&��JK{��U@n��/	#�HY��D��#n��}_��ޛ��?X*�����!�ҫ�I�I�,i_\w���iƆ�*ڂ�"�}�695L�~��J�x���v>Κ�5s�4r�׎0��7Ԓ�{[}nT��r0���H�1��15����@�ub�!L]�����r�YY����>BEoم� !��00hf ��~������髗�he5���lde�K)x��C��yf�2T��:N�~޷`���8�5���uK�l�����26�=`5m�(ζ�)�q�Hht�dl<��(�w�B�L?�wQ��@����B�%i�R���B�IӆR������02Â����8��%5s����	n1$���#��PBr���v��p:�
x���I9��Nݭ<��}b�|�*�����ڮP��2�o�������_�%���+�>2�^/����h��%�`
-*C�7S��q$ѫ�5R��K�枖-�[U�8�Ϡv҇���L/�z�-"h^�ph	IG}�u����lz66<%��Ϛ]���X����TO+��5���57F�F"l-�*#3�Oʨo��|f�A_H��"�SbP�_).o�m���Ǿ�@xLW`�ю���Q�����S�f��$��b��<�c]j�Ӱ��_���*:�N�O�;�:h.ԅ�kQY���$�.ari$zO�7L{<bF|0�@y1�N`Q�}D��IYY�	s7K��as���A�z��Y�<!�=yi`���3�5K	�K��Eu0���B�7���I������c���-��5�-����N+z%/��da������W>��W\�i��ҾI�K/Azw�EU�W%�����l�������i��ӲeE��`D����GŻ)���B��	t�aY�����4���o>&!7Fn��g��$��F��A|S�!�1g'�ԚEO�k'�g|�9x��p�����in�OI��p@:�[
�D�/�V=\����a�UI���ȳH$��)�EA�Q�"s�ߎ��Ǆ׎BX�9��Q�GIP�M�󊲶���"���D�貃x�;���u�-��y9N/R��i�v۹M��唃4VF���6�!֢97��<e#�>lO7�(�����t�֦?)��P����S���ڳ( Òs,�Q����$cKI~Xr�����*��J�fee!@��9"U�9p�S"�$.��q�T�Ȓ �^X}�=��4y�!��XHㅬ�:]4��2�漗9����0�討�������=b87���U�V8J���G몰��^w�<Xx^71��ɞ$nmr�=s����$sʐΩ�E,e=���F���Js�l�^��1�G�/���gR�ܯ��k{dUOz�eD �RIm!3���Z�6��P)�!kڤ�>�i�K��G��O)t�X�[���߻�(L��OL�:���3y����p� ����
���n(��:��po��J{�|m,���>�l��M�B�q�~<��`ߐ���t��1�x��8q�o{H��a��A����C�l�f[ w�%��tpMh��x�?���vW��T;D�ɏ8��Q�e�ԚiZ-.:
iC��/Ҳ~���v��� �L"K�v�7sU������^�gd�g	�1]�<&��ܤ�/%�6W�[2�~��{$���l��D�M-��P�e����ŗs�����x�'�J���lB-�^	*϶@�j��pO�0A��p����LS��R���f������y8��W�~(�w�+i2%qSIЌsu�v���� ��K��T�����#�e/;���l)0�2���}������.` g���2(�>/y�y\�/)J��j �	"��� ���>/�	;�J�(QS8=�<�5@��k<dgk��t�֣rY�����"_��>�HSER���!���q�F������D�ƍӧQ�cSU	��Ȗr#e[���Bu<;�GOZ�Y3��vhju�l�sN�?��Cn��3��L�]P��-���O0	����]�V�h�8?C@��������qX&p#�!+@a2�E%m�W��F����*��Fv5e: �OgD��A[���3�<�E�]��۶��VK��U��z�4FJ�&������{.�����lŎ�ԃ��Ko��8�^[�8.�h���|{�q���-ăj�v&G��Z���W�af���1""`>����=6geG���{Ӧ{�c��k�u�v�Sk�7��Ac��HQ���L#Am�G*�B��ïx�T��Ӷ��o)�����Q2��H(��"�<Y�Hb�%i�La^s?!Y�Ԇ�� �����= ��W}|��u�\��?�#^V�����uT��\�q"��{���ը�I �:���k��:0e�H�-2ʚ�)֥�����_���l���[�0��gl�<����įU,U�[�~S���ZDN�ALs\�C�v�a��K}��c�p�e�n2����h�p1�"����/+���l�:�eAxtN�g�D^��R����W��A��� �;� w�������P�2�B}w����K�9�e�\Cҥ�t�*�Z?I��ǧ�tR�-H)2g^Ϛ� )&\�����"���XQr�U�G�>.%{g	;��ͼ��a�`���M��b�i��]�纔��şĦo�����!u齲����j��R�ꗐ9'�j���¯>|�B�9��]w��aJpRV$��n߃Ioqa>\�]+����lq�\������ �+~'�p�}� Ӿ�D�=��Ӄ���������ƹ��g�Z<����)wH��
k;�n]����k�>�
�HJ�2��U7k��">7+���Q�߮�Q��%$@rL�X8y/��$����M��2>�Vl!9`��׻���h�@��O��x������.�=�G�׽Ӓ�}q;�-��np����i�گ������,�)w��Hy�kQ�Y:����I��/���c��F�����<o򒇹m�T�ʾ(�~�|��Ε�Y�AN<�g �V��B��F�z�~<��*ϵV�����h,F��K ,WrM��;�|2K8�;�{���:M*�gq���b���ooo���%L���J�]ĳy���v�����O��"ӑ���5��rb[�hJ�Mck��s�s��y����������1�
Sӯ8�2p�����.�t*Ξ�g�JzC4/?��I�nz	.
��NԪW�3�p����sƧ�:��H��D�j}m�Zc����~��x0%E�gp��~NS{V����zQks[`~�^�kI��ݲ��K���3��sU�!!w#�̜C�i胐;v��]�xѦ�������]��y��Z��g��^[r�	v��a�w�I`n0���\�0��*�-
�`9$�ޅ	8y�niu��ɇ�0�e)z�ou��X=؄��'!��B��Q{��V��k��$�t���r7�I�ʻſ�k�C�~mӹU������z�jQq�=&��+��o��Z3���\�*&I�K�ɚ�.^!�ך}�� 7����*��I-�~D�yDٗ����o���'���ݘC��.K�����%h����fW=�#������P��O[��L#[��!�vA����@�S��Pc<�oY�F=df��Jɢ;�:�$T]2�ݤ�U����y9∀���$,�U���_\,��z��,,�$#�y����Ɵ�������.�q��OH����4�1�^{�4e���Zq�x+�Z�1��I�x�N��>Ћ>I�\�R����F��T��X�?�+�ۨu�M�F^Y4!@D�^��ʾ5��ejP�1�}.��X<��Y�\�v���h�V���<����c�9���%i���p�H��{X�h�pf���J�l���2��b�Z�Y�h��R�C��a��h���c���\�jI�K���m52s���_oz ��l�o��>5�7�y����粱��n$AQ��H�;��t��Km��.��'�nj&"(��#��$Y�I�c&iCt����!@W}9���)�z,?�X�&��KT8�y��x"�I�a�F#&TN*� ���cZE�E�u��&A�Q�(�P�z2i�D��K)N���Q
�r'V�n��Z6����H�w/����m)���q��p&cļ�A�Ժ�+}QJtQ	%�fCQ%Lx)�I�B�N4����K��!�?�Y[d����=Qu�*-���r,n�\������aCmU>t�]KI�8�����Z���r"K�p���u�o�g��_����jS�[��_���e�%<k�A�F�= ��D�6���6ƻ?\��������{&���;K�72*�
�pH^�p�;�H���i�S1RK�D��m=s��g�;p�=O�ӽ���E<��M�(���v��W"6�Ȕ�~N[@��Q�Iy;]�IT�
�*^�㎵�&���Nf�d��]F�{ G� KK��L��^0s�1�y7uf�'r���r���ػ�����iL^���#��̕��<F5��u��*Dz��b��	��i�p�H�;OY�L���!h���������#O9>u���~�-a*�K#�L���}�� �-¿�[�өt.�pE�D���&,�K����a8�+���5J%N�~Z�#杭`B��I����/�tCM[��W(LB���!��G��yT��J�R�X��������
gY����+���aɸ|�Rp3�� ��QU'8�x��9P����F틪��m'Oo�l	"�<���wH�5�>��`D"�����V�ˏ�{��ٝ�M��u�n��`�|�h\�n�ȣ�� �b@����g=0������շ��v��>��kD�G��sɅ���!k�sA4����.t��@l�<�V	�J�ϋ-zX�)%Ð@k� O\`@�˾����ݞ����mf��[l�en���g`�'��p1���ܘ!ک)�K���H$n�#���$��F��A����.�َ$��qXRp�<��t�N3�	�RK�̋�h�8l���k�EM]�"C�[�ȷL��q�Hl��k�A��D�FZ�_==�yf�}�Tt�����Ҷ�$�K��p���Z7�ITY�5���-1-Ƅ��-�xj&�≟��/��Ka�K����i2�-�y������!�MR����P�̏<���gu,d�x�BK���}őe+�c��!�u}�o��5�ohL�'�3�+rw�ݼ{�zn:q>�+Zl�T}i"�+��Y��Vx�u&'�xt��t�5�-<�[5&��F�[�Ӯ�X	�Ѵ%CEQY��fk,�/�=	,d��W�"@˔+4��<i8�Y�+�rK���6x�k7Y#�rY4-û��������-Y� �UgS������U'�[d��Nu1�(ӳT${�����
�i�|�@Är�;W
�jRп�a�~�E�+�0�:�gV-��5�5��7>��Y�DDԽ=H.�����֖٢��}�Ѹ���C�A��c_+������^��v�m���^6W�x"Ƹ��u��e�y��>�@FU�yi����<�I����IF �fV��)�	gӓ吱��z7L�?���A8wЎ���. �\3Y���H7 Y�p+#�n�nJ  $������u�������8��A���=!N$�~���� ������8x?GH�Y� ���M�*}Q����em#��B�8�	�@�-FV&rZ��;s�n8�*���"����^𿛓�Ѻx�rr�������2��y�m\=�&�A�1��KOn�0q9نօ�]gr�^�v�2�*�	MM�Bc�+�;o�JX�A��ȋ+E�?E����~����Ҿir*|ߪ`�NVH�M~���Q>1�?K��d%S�W�p�k(�ёs��t��V�T��'MzI���q���v�-��"�����#��Y��姏��ܣ���؁S�-��S��*���P掀ѱM�j�Rv<�$�����fY61�U ��=�gC��5�2j�D5{]�!�QP�bkױ�1�9��	����7��J��ݻ|�芘������2�*Se��)�T���^l ��6V��
�h3���T�K��j��k��qh�Q��,6w&��*���{:��� [�jKoh�/?<N
KeJ��qV]�Bp�Ӭ!���(���ʀ�4x�;Bp�X����V�r.�Dx�8�Y�bX\O��x4�Ő�LB�-`l�����[��(v�^�ky�&&��!��RC�x���۽O�>�������e�������Z�m���=�?�/OV�nz�q�,���������u4�9jz&���� ��E�<��xE��M���.?qT|N��Ft�
��Þ���Vm�.�1�la�{:M��n�ʲ:~2����t�$�r�;m�4NV���a�����:��Y�`�ל���<Fw�o��%��n�><,�@�U^�'l�Lm6A�ne����oY��*�q�0d���4sX�C\�.Ծ1^���e������b�uWI��CM	��n4�"D�^[m� >�%,���Z�������͞2a2#��7h�B4곡���X�����1�_��0[��gz��LG#�1���%C��e�'�O�@�SQ����`��!�q�\�/�oe$V6�������5�/R��Z���RM�AB�unsHE\��xd���H8�r��W)y��$9GdI�����7g. �whj�ި!s|{�k��7o-�#�����?������ߦw��%�K�:���3qdTtA�IK�~J��T����0�X�S{C��ǘ�c���վ	R�x1@�k�pr2�I@D���O"B��K��@�``⧒4Q�E��F�:���s��M��CT�qC$l�e��/�]���3t0���-;Os�yQ6b}��'��As���e?��(c#�;t�$:bZI����)Md�-ss�y����+~ v��^���G�y���ƛDg��<�v+_�����L��N��������'/�I9��qT�0���H�:kQ"�	�=F����J��#��V]����0'��C�ύD���jf����֝�����嚐c{���l��5F�A������(� ;�xR��S��(a����Cu0s�;*`��n��� ��O�T�!U���a#��}9���S��LCU[�����1\���;`q���C�x��)k5����Ba�aƧV��aJ����|1�&c�UZ����C�:$�yѺÊ ���Χ�V�1�Y@-�%iM.�`/��u
/c���I���O�h�^!"F��`=1v�&}YW6]:|b�ű��?��3�+�����E��w�����I���Y��ψ��g�xu��Qb�=B5�h�RM2��W��/����BC=Zo��Qf86�s�B��7���*Y��b��t�T�kq�4��Mk�#����>I�kU�Yߧ?ù�˧LL�"�����oꪥ��Xڣ�,i�#�fN��U���h��k�ă��8E;}}�2N՜6C�Yn1��e�9�4h�,����j�L�����Z
?����a�}�,�_bA:{+v�9A�8
�Z!2�L]��&G��{�{D���n����y�;��-,S���zV$.�d�D�Ч0���^�PP;�p��}�f^P��[1�|���R_��%�6<ECq	��=�2�xh��o�R��0Z8�}�8��.���Uy�;u%��	�{4����� �ֶM��}+2�
��ѐ$p�3k[�d �H|�R�{xѭ��K�8^���Vx��*�U7#�ʙ�����ߕ&���/�������@֐�,t�Rfzm�9M���#,\Ո3��4��� �x�r����ZC���Jx��ң"i�w{��2��r-��=l��o�t���?��������V����f�APC�N�i�M?�����4��f�=x}.��t�z�I��ӊ�X$q�?c�[�L�Ft��b��@�+��������!�=I�e�b�0����x30m&������u#��w�W(�v������^ꚳNގϐ�+
�w& ��ZD�笂��J�b��1K�
K@ɰ:� ��e����Y����,��pt@������ܤ��>oh����������@��5�i��7�j�3��)��.ء��t�&���}X퀆\�Z�tl�� N��gᚻK�rJMӿ7L�����o"+f
P�����M�[9>MV�?%$G�չ������b3��#'
{���	��_�D��T�r�a14b1[6�}9�
OY�]�jg�k<z��U�y�kD~�������!j�kʪ�r��z�P�2�C��S7� f�G�I󌔯�N_GT�Nn�ˇ%�s�C��~	 ��?|aU�1�a�yL7����'���G�
�i�|���@4�����]��n���x�M��䭳@6��l hs�WQR;i���Ė���8�<����]L�&눱a7�/��,z��J��ƳD��^���w��di}�jXQFOY+)�,yֿS�B���6�^G�cr`���ɇ(�S�@d�*��H�Y��p�����-��a��<~���Gr/�5��nC
�"�`]z��KHFK��\��Ɲ�
��k��躢�rZh��*N:�[���x`2�Q���+\}xb�V�a��cޜ��������y	�\���n��L�k}��Ҁ�n���RG[9��y��(@]�Ql��&�����<}v�;WY:Ix�9Š��`0a}IO��i�|<s��5�Љh;Y���N�_���[�g�2F5���{U(���Z�WER�e�+�Զ	��#�0��PF-p�i�;��;1�	B{]Q;��n�)[�)&��hbh�İK}���C��/KM��9��/�Zq��Ƥyޔ3�6=��ܢ��Y�56��$���������� ��`,����
J����c�Ɲy�bw���}I���>g����U,;sf����P[��D�%ƽ& ��T�_G3b�6��u�=Nv$�Y]��{����Ux���� <;=b��N-Al=*/9 y�;�+"��p�|�^��`�yt5�(;�8�4rv�+�.u�R�m�7d&�[{$3��S���~�a)��2uc��D4o�%�J���&��a��^B�n9�A���%`c��m�JŹ�2$s��Xރ�JӮ��f#�]u��V�MJ��.��0�F��ωu/B��ם�:�w���8h��M�%2���<}.+�c��#=-�W�v��K^J)ĩ�Ҡt�b���j���b��'�#����J��)�t�@'���[n���F�>�y>�]�(!24hv�� E�x6�_F�Ϙo�x�Ϳ���P@O{)xE�a��	N�ӫ�O���:tԡ�3��؁��~>4J+��	����촘9�j@�>ޢ֟�d�D�8�$�}���^|�&���KRI��Ym���p=��1��|:.1t?@��k2 ���<a��m-jmG��w2ڦ�!bjM2���ĪPŸ�ҷO��9�U3��m�� ~�Pg�g����k��ih��f�/��ZԚg�Dl
�¯�Xpz�����8咖Y�]ٷO˽f��/�Ȃ��-�B��Ȋ��an�9)�����~2�C@W��� s��}�}�r�U���l��N��J�/�;5�_�⍯�f������߳*,
O�Lh��'.��`Pi�>��'�w�.�����|[F�!oE��(�
\y��˨ڙ���7&���MW���l4���ۿ�Q��[��c�0ڔ �9,�G�ըp�3�#˸�|�:H�˂������P�S��,E���
�~�ɱc�u?�b_,�b��glB�l����@Oq�f�i-�� ���j1��/&$mQ�2ɾx
��VS��-b_�J�ŽS�<���\��Nr>wj[y$֊sYR�JlWE6"��P���1e�iwe��Y��֗\g����LB���f�*-�y��ϔ�mN�n��.�w6�����z\L��#-��Gҁn�Ǌ-��=Y���n<m���Yp�g������&."�j���pc�@���.Ͽ��4�Y'~ӻ���V���P�+�'� �*y��C���	�����Ѫ/D�\2΋�u��Q�K1<�'s
����E׳���wM�j��'��i�3%Â�y� _�������<��\��7���q�. �E;�`����4��(������`��׆R�����-o��6~�Ў��)jC��g�Z���]���WБQ�}!P(Ho�u��(R�nb���;��(�������F��V�$�QY`h�����64�	��[J��!�'ױ&�=�s\oOwo��(\�)��b�\ƏA�%(vN��g ����3��]�n�d��5j��od��;쬆��%�Frl]��N�xx�Qa%?Xg&_�(�vG��됱?�����P���]!y��P6�lጃT��4�Rօ�ѫ�]�,̋���:�j���
�dԊ��6��l�K|d���&j$��rҁ�N3���phZ��ɐ�8p����X�#�i���=g�QǤNwH���(�<�k(D��i^ ���f�:�����:<����*�(MQ��#����V4�{r.]\�ZoOp�����<U�c��3��dm�`B̋Ӭ��\��5����GR#�rg'�`u�Cak���-f.�?ĢU�u�uFY�9Sҙ����'�,�F�@��Qi�K�rm��l��{�;V��@L�b��Y�]ש�*��!���z�&�B�ڰ��lp��|Rs��� ql�@0H>��(ֹ9�t��{6�5{Ѳo�n�l���rr�����T���r��%���= &0��b�/�͏��қ�ӭV(�tq ���Rk�`
�@��E^:O\��F�1l����M����H`"fR+�q��1��P���V��Z����~�s�:�0���sB��ٴ�,��f@���=���EpO�u��r���3�e��+@��%��8��� �{p+崕�p�$PG�k��Y!�7��dla��K=��J��Cx���������r�1���������ar���ʴ��w���y�ӟ_��	8���V��E�� �h��Ho�)g1�F$�|ǀ����KW��.�u�N]����\�2��b�?q��m�c)�f��'0�ΏA�bT���EN��]<�9A�3=�_���y��
���kS�v���Ը- ��O�h�r1�w�"$A�P4���޲�k����C��_�ɕ1��L�-�����|T��c��
�)I
��ʣa��p�t���݀��%G,j6pG/�ž���_���rѭ���^~�r�.tb#�iP�@ႌ��>	��h3R#}V�t�	�T���ǮM���"��ld�*�{r�$�i3ևv
���/ρ�|�aχ?�EB*f����r �gW�ǫ�8�x���[��<,� ��A���qX�*�!����2{+�x���6.jJ����4trZ��;�SwOQ�6I�a��cțP3	/�Q��Vt�)k�ڙ��֢�d+�M�*�|<�{ 
���B2�bjO{5Qx9�H���<���,)�z�'~JO���`v��ڙ�J;��8����� (e�j#�;#�)t5J�P��FHgz�Xg}��TP>�4�ދ*W���Z$X�Fx�;��,}>҅����ChL���PW��8����*����bٚa�rt8O��#��C�=xj/v�Z[ě��R�I<D'�5�3�)9F2��tt��m1�A��3����@�e�q0�ݝ�������{��xOYۀ� }-!!쎍1>0��{���7�z� R�=d�4t�?���h�`uת�j�I"LW�?[a������2���dn�|����g���J�[%w-�5�Z<<�-g@��ɓY�Y��c�+��P�����ђc�m|h��Ў�ٞ���|:h��6:(V'�x�q�a��&��0d�9�5��녂]�!��!}�$�=Z���Ҳ�!l�
�Sڳ��6���q��1[�}�4��UR�|��?ɵ����eDj!�U�O��:y�3yL
�e��Y��qs��EE���x>��.��c�_%��$O����O��e��s�Q���Hv�[��*C^Ұ8q�M��`�e���V4[�]���h2�#V��ͪFʎ��?������F�G:UsO�4�Zr��urV�`��%686Am�P����ܳ��M/n�?�IO�����ʬH�'x�}-6���,$��]֭{X _Ʈ̐0d�@y[�}�\��x�I��9f��kPha��C����x`�,>eT���_�(�	���$�6��������H��>|2m�p��*_P��V�v	ӱ�y���p�~۩t��8����r�b�jb|�髆���ٵ�����2�?R�TX-�*��'��.����L��O�� @�w2��]^!�ʮ������h�ww'�g��{��(EľL酹�?����
R-	����)���>�̿f���>���_$�p��i����B3;�0��Z� �o�c��dBѺ,׹��L���Z�p� ��l���8��:C�m1$��W,�f/Ν�9�IK���0}������J���bn�y�@���b�����/�<r�����u]Q%�*��,6�ݙ��w�������2�8p��t�9�A5�E��v=��i#��"b
��*/�TgĦ�s&ſ�^Eo�:��'�m�$��kFxIt}����U��&���:Ǧ�27�D��z:���&���~��~�z��S7\bӬ+h՞�Kj&���v�ɛ���}v�^P�C)c��wA�7P@	�G�$�j6��h:��N9�|!�j}���`��w���鹞����#�N1�|P\�?��ja�A=�X�i�A&'�jO���SR��2���u�3�*\�����o<Ds��pg&�v����nzҹ�\(�鹱�h4�ݍ�0�U,m@�3_��t�W}�\D����v���lr�T͌����K>�ie���mܱG2&�7j<5i8��<N��<['GNy�A=Z��K0-`�A��଱kĞj��v��~�k��l�Lp�sV[�j��/�5T^*����_/��=�6פ~h��h�.~�|��+o5� 7�GG�q�Jװ��T���'���9G&�]�]5lHtߗ�\+\r���dw�-�����E���uipEn��ws}�B������\�w���n�sj-,�&���c~��r���o��E��Z�$���4��-��f¤��U���p���s�akaZ���6ǩ��WI�VS���5C���O�i"�S��n'���>�T䇬�D�,t��naQ���O�Ӿ���ԋ�G� 
oy*����S����2�vNP2���Q�_)!��ok�F[V3��%ԉ����.���ۚl��Ҽ:��w-��wg�]�0� �"��N����Q�:�4aA��4<�q�8~0����+�vM����mX@�̄.��ƾ~����(�JsY�*K��O(aKw�^�� ��!#{ë}��*7G�!��n�G���5���S�����ǥԒ"_Q/�:�k]�'"���Q�4�x<IB2�e�gd�j�_�I"f���$�]���
ÊL�}V5M���%4q#�	��vg��-�=4�~Q�
4��X�8/86�x�Nk��w	λ��[[�f/����E��H�-~9V\`���|�#߬�� �z�,������<7�?;�v0a伙j��b�RL(�7N��Ӆu��
Цz��ó]/6~H�B�EncT���Xb���Yd]�����Y�~Lx(pT�6��(�eq��At�Y�=�d������(�\�$8k��<T#���Z�������g��J@�>ˤf�������A�mzIR�AE����%KB�N�"$���:eǉ�E��%�-m�l��{Qȍ���l)�d�DԈ��l�
���� \nDf�߼��Z�n���\���5��8"~��a0G�;q�/���x��o~IW�ץF�H��"�n��u.?(������O��bz<l��H��#�p��=t=�Id*�,��O�w� )a.�X�Ӽ,&ED��GL���զ�?��F��D�'g"�Y��_�5;
��{}����$K��I�n
O2W�L�	��3��8�`7۹0�#��0�]��0���]�I܁	�D�0"MّBz����|�����*ᇫO1]��7Z��3�B�j�VF&�Bv�����h�mr-w]�J��f�@"9��1���vu�]q�q�P��B�xQP�MNs�P��b�� �J��<�l��<�����z����&B$��S�Q��N�8e�=3�ۜ[^Q��/`��L�A G�f-�*,�U��M/�X���2%L��{���{/��i�|-X��D9 o�k&U�r1���,k�QghF�Z�k��C�?4SķŹ`�\�.N���52����2�B�����G pl�R5�*>�1�� )&�q&M!�/ui�˖ro\�d4������MlL�'�޺=M+��g��Ip�6�p�L�J���>�F�~D{�\\�:�P.C�"k�u����dJ���y�Rv�
vw?t�vo��Q��`ƠF'�,n�}f������'��XU��f��'�x0�I�W��6E�׸�4K��p�@�Oń+ℰ~:`��`×� �|��}yY]L����֏��&a�w��{�� �tPW(���z��kxV���ʣi<���=�6�=��=�CNy�!B���AK9X����@R�<Zr�8I}�+��,3�]�G������?�NT�U�dR��}nA�����t�݆���*p�퓖��F�eiQ�
�PX.�u�
T��$������G��-,
m�B?ح%���ǠԞ����5��@�����. i�(@�h�y^#w��o�,h姶��^����R|�y���x�#FX�fh�j�;��gV⮑Z���(|C��N�Ͳ�kǜ��0\���-�4,��G���[ὅ�/���謔ǽS�2�5m��I���#ƩP��5�N&n� ?"6+�iQ#G�r��o\:������޼�d}dK�8޸)�yB?͂?�W�����p&L9]K�p;������F�u�"X�t���(���9L�ȅ}���QW�A"]�vz:E�ّ���v���݈rF5.\H �,�g��rJ�ʺ�����#3�$�b��(Z�>iz���V��Yc+���o�m���u�Z!]#��m,�>�������P�,�5���b���+���܌֊W� 6�>�@�g����A�R�:�\�ɉc��퍆}�0b"�>�P��'����cq+k[�k�� �ޓ��ai!��.2.���Y�b��+���.��'��y�`¨ �!��9�xMq��O�vȞ���56�@���M�,��]՘�Ij $#�?q!(�J����o֏�_H�g(.�Yl��\����o㤃Ky޹�V���1x:N�F�˽G݃�ʲ��yW*����j�4�V�]Vh�_��N���#@�CB��X�R%,�d��C96[��L��@b�9�W�����skZҴpN4g6��W�ۄ�OB�-"��ta�a9��T	�%�7g\Ꮜ��"�D�8�4#�Jh<v�?��iO�q��Hߐdĸ���e7���x(M "�������e�q�Whj�/��G���ćyd�!����Һ���y�i�mE�nW�&hg{/���zG׋�P�J���5�;�t���꣬�z�4i<x(%����:2��Ѫc��{�cL�ݥ��'�;���|�]mu+�*THf]6`6�ʝ�<
���b�V�+-��,
�< ��rr�s"���/�8xb���~A�� m2���!�7��m�}�6G�$6o��h���+��~H�ڽ��f��d	�R�!���x�nI�9�W���dv�g�ʿ�7��gUp+r��
�[�>#�f`x(Կ���2�[�H�g�&0�����Qpx��_�㿲0��V�R�e��\��=O�Н��d�H�U�g�����}���*7�p�%�Ժ>��JԔbQ�J���+��V-�0n@͚`�LL���Ū��fj�������<N�mzx{"�� ��z���s������G=+�\��LC���)����0P����lh������N�1��xLz;�R�-[��L(5�O!_���C��0��*���4���	(�R�W���22��V���42�q	()m�"9��R�����O(�ƠuԙސӋ��#��fD\P�	��j?O���6&ʹ��tC
X�g��íy.��d�I������yshΖ�N|�C�t��1�Jk�?J�#����`��=��-��D�J"㌙�p!�w-�o�1����b�U�����"ƽGN��7����^��w ���LL�ր�ƃ�M�^�#<���Yq��Ľ���Zt�!��L&�� i��:��e��?�$�f���&�* � �:k�I�$��ε�(.��93��4��M�,��kH�%��پ��|Tc�g��r��+.#1�GLͽ���`d�S��F������}0mX-������xg�]�.�iw�'T�q�ܕ5�2T�4����,,>��U�c�.�j"w�N�e�7'EH����x�+��s�ΐ����R��1�jQg:�.�M"@':��k7�\�	�%/̈́}lbx�y���~�QI�8���X��3���a�����~���,�e[E濍L)��{��@���X�)�e�G6�?a�NNo��|���Y��RH�.��?tQPXq�rX�}��$��5��d�}L��)=��){�R�k�!#��Uuj�Px��
��1<;0|	w��8�}fh��GpV0���(��;/�C"1�2��Uy�O6�G�Ɩ\�Īн���9+c����ɼ���8h��QIk63���7���[Ō$j�}֌A��"�@y�,��է1�KU�9�������V�ɍ�cs��TM����G�=ǂ���f��R-Ѵ����v�x���e�靽P��&�B>�䁇*1��36���x[n+��ٓ��B��c�B):5��7�=+ܽz�?θ�a�$�^Q#.u�3��i�������D�K�?��ѹ���50��34��D�W87��!�]���y:���4�:Q�p~��2���5�/��&Y��Y�z|As��m<�<��� /�8��>5�����cv�U���i��}f����N���%���x���mV�اn�&p�{�W�栣��	��xc��8�uX���E��h��6z�Kd�7��?�B~�P��Q~.hD��s�-�wOK0��7�}o\�,��@�ݛ��:eND�DUt��J��4��lQz]��9��GD�))�"V��Ub�l�ċ�Q�Y0�����{䛑L��I�S ��sס�@۽k��Yķ�ʤ����A�(v�-ft�N^�CƆ� ����2"4t�xT����3��z�V
ؗ�:Q��_�X�r1`Ȥ~��e� @&s�.��>"��xD\(P��\�f����Q~Ft��؎��|U��\M-V�{�|=
�;4J����Bs��㠺��~X'�Bj���?6>���0����#kd�(�T�5��1��z������nX��|�pU*��nId7�]%*%�	�s03(ޣ��d�ᒠ^`�ی����ZC	���Tl��B��h��Tx	���ޮ6̓zWR��1LO�h$�[�t26d�À�+@f�D��j�F!����% V�9� |��	w�L=�ȶM��Ջ�k�LJR}<���oY;��r�3Upؓ��w��4k9C$�Q~y��"����y[V��r�;�UK��Ŗ>��k�����;��bUn��Fߔ^�`�j�F���UѦ�Ց�3�����x� ����i̓[D;��H�<�IfF�GKC�)6(f����Y���7�K+$����'����GL;�m����*!Qo�'���槫 �hG�����&�Lw����Q��r��h�<Պe�|�7��A����)G��N)r��GH� ���a_gV� ���mFH�y�o�I����uK�(�aؾ�)⚠�<J�%Ơa��q)��\g-��.��@��ptKI�Oz^"+��j@����Ã�W]�#|��@�*���z�nJO�d�N�[��σ�hڻy~~�����t���� R,J�o_�+O�wS �r?��Eo���bX��d#<��p'LGW�tLGy�^���3�bv�Y��iEJm3�ڌ��Z��|.>
�ݰ�*݊5�PQܺ͟h�a���jO�GF$����0ʁ�{c�ز����/;�mNw6:�㎵�m�����J��N�~4��a����%�Ǭ�qA�o#�4�gA9�� w1C>��X������g��6�gD+��45��(C�������e��*`�;��Lq:uP��T�%�q2*.A�X���Ntb���a>yـ��5n��7]��d�\ fPv�H %� ������"��R���;�,4/�Q�A �ϊ�� �)��.V>P��C�U�E������g��?߈���U;g�ͺ�h�bǞ��������]a�.�;v�?�a�u���R�p�w5�ϱM�6��&�!��'�1�~�V[p|�n�zx~� .�T�DK�_�����L�����;�bE��Q���-�q۸Xq(DZ��G��Ѹ�ݵ]F��i`X)�$S�7�}&1HV�ci�G�`�ӁpQ������woӌ�r_S;TX!���! q�ǀ���o[�bG��Kq'HB�2���~)@�����d�
i�e_k��}�DW�}ɔE	a>I)W�)�P ��ʦ<5������|;�3�#�y��8�r����i;���� |��@�[֟��D���Y'3��$�� ՚L�5��͍ܝ��W@��ș���Њ����e\a�uC���Ƞ�����"��~��.T���	ܑ�6:�L�,��e(���p;���b�t�F���D��Y�i:��[7 +p��d7���*m߫�-��	��p2iRx_L���S��x��kb~mg�0�1��0��YH�'@������^�p�z�G�8I~�n+���Dٮ�hrx���9����բ4%"��|�n?��)n)o��sM�S�,ؾwDk�C�6沓���v��G��)���R�Y2n!$x_���ύ(ڝYY�u��e!��r����Q��[�h9u����Yq�� v2r
�$��N���.p��`���I��l��bX?O��ә���'}g�!�6M|�&?���JC�m�h\>���FS)�b3��d A UJS���ټ�,�훒m�� �?^w�v�x�7����+Yi�tC�\ʚ��������Uo�
�N�F� o�H+i���&i�g-r��Gs�gVt��@E����erHJnt����:����~��uߚ/
�5�&���\7V<­�R��8�P�#�;����SF'm�d�90@���(�Y��ME�&�����h�i˗��uN�n�c�����*�A7rgԘ<~=ۼ�'�\�ai��:�3z���)��ݪ��K�Z�8�����G�rAX�ܦA����؝*�Ż��,���>�:@�Y�*�Z�gNi��hmK�ީ^�m�*�c���))����u
0��"�l]���P�ߍ����@�#\�*ӷAZ�Q%�X^	ñn�  ��sR�������;�5kY����}�N`�� ?������	�JS�y�~�pO@�h>�,�=l�$�{c�dDN��A�6�������'���D�b�֪
;[G�x�}))�j��a�i�U�/*���A"gu4����.Xk�6�.&s=Ei�ٟ�`�|�=��ⱌ��'7�H-�t̥���`�K���R=�R��0X��k?v��\�щysqi||���@��y���L�ݤ��'~���|dA�`c�6y=�l�[;���b����)C�ؼZ��&�4V��$��ZH#�(����r�WzY��[�{��Ty�P	?��0��c�SePߎ�%�%��_i*.��<�
+�7�9���Ui���T���"�1�N9���7�9h�9V�.����C^3�D�N.�쥕!�X�E��	aP��BK��_e1�r�+�:kH���h{�cU�b����/��
e9G:�,S�E��A�-\��Z���1N쯗�1�$�
15��1��"kvL]��q�@Kq�@�q��m��m�Q<ڔ�7��D��>�i�}}���s�m�~P}]���rK|���`=�9
y��K*���h\�Pn��Qb�iU%�2#����|�V�����%1���D��.8�P3�D]�+��}&~�8K��9��͡,;T�!���\�Md�]�BK;��7K��WS�J���G��&�y��� ���������s�2�$yZǴ���\iE����(R3~.��Кx�y����Y��KތL�7��"����K wyV6Őr�N�a�b�=����_$�y��R)��
�0U9X
e�5�W�����(�1GX�,7w��e"A}�_V��A�s��5sZ�����AC��o[܌To�Yb6*?@�pl�*&\��!]��`��_�=������m������W�#�	4���$N�x>��T:3W������qt�M�*��H���N��'\����ȳ�����s�q�!+`��鍓�5q-���A���J�Ṗ��YO�A_��)��u�g\@����PS��Ś ���7�*�]��[��+�3��Sf1A��&��M��&�������R�q3�j��~�5�euz\r0�)�"2�;οpM��)�Qγ�[���=����8�#+G��R{���Sa��J�Kiv�ʳ�����I��6�d�h������'~��AFꓐj9�%�R����3����ɑ�Q(�\�A���^���^�ά���Gf�����:�(�si;to̧m­p<F�D Z�ehe�#q�X2�{�����ڊ��Rϻ�X%4�,�����k��oIR���Y�b���_��X\���� V~���[7�G+����D����%�c��?W$[�a�qGp�U1�%���|��_q�˕LҨ�hT����6�q�)��V-��� ���1$�BǏv�P0ψT�5 !3��]�h(�N���j�ZC;���*
^u �ы�x��e�b^�~b�_�!�~��,^:��QO��픽C�cَLao���'��j,�)2|��a�e�렰�ͦ��}D�_�f�h����mOƽ|�;�h���fy���i����-i}��FЉ�b���O�#s�����5��_�Ǎ<�*�`���9o8{�^�j?m�#�}-^o_�X��%��^���{""�`8���$+�Sj�h��S�X�T���V)�������Nm\��=�R�o��!H��_)E���6k�`R�NG��R�P0@+9��PJNqv�w�<o�����>L�Vz,\S5q���>�֤��SZJ�d�RL�kϡ	�WҞS�p9�^��?y����`a$�B��mXDY�x�Y���|\��g�ɉ��WX��[���ꈺݘ�-S-)��Ə1��,-��kB@�=�7���c��Ņ��k$r]R&��M?KU�xb� J��?�TA,�<r��_Ā�E����apy��� ��l_�%��1����z1IJn����Uf�rH�`�ot?~J�ˌ�o|�IfWhZ�����O5��o����� ݁�c����y�[s�Ҕ�D�`�
ӱG1$�-���M���I��?EA�4���?ؿd~�����z�zB|�q��z�&�GmG���{�19��L۳{�y����`K�
���v�-=����j����]�p��sǗpO��0��]�����N�:�=~������%���i���R��Z������~�h�W��,����E ��������8{�4��v�G���9�������Ĭ׈�P����>df�>*�no!��َ �����d�Z�$��ьj
��#%�CRʈ��W��%6��zej/gif>ܳ^�U����TJ���	
����l$���
aa7X�H)x����Ђ�_3Ų�����8&J-s䦜{=�� T���z^��~�ה��Y_�ݺ���p���t��E�#U���;�q���T���Uw�EZ�����%���p�iʖjo��ݏ�p�8q�����YD�0�5"K�b�ww�P|X,F�4��L�k=gӥp��j��o���K'�el(H!S�/��]d�C�������l����N0��+�1/l�M=��%�����xص���H��z8 4g����$|u�R�������Պ�*���EXI
}��Z�E�=���^C����b�����bԱ�)Q��prΐ�G+���Q�9Z�m��T��:r��G�d<�l�T��b�N�hL�@\�|}���;L���w���,�+��/V�(� �h������s�_3�Xs����\!�~���h�ΰ��N��\�#�8+BR�*��&��J�S_6��w-0�F=������E�&+磭-�7Z\&m�F���I��x)��#����M�s��`���.4����O�r�}����mɺ���j�]�!wR�6&�mû�:~�X��~�6��;�,�=��plp�������+�����������b;s�0�݋X�oN��=��b	o�<�Q�B�L��N���d�C>���/v
8l���jﰽ�r�S0��8Qj���T�i2}zDD0� |�o�'��F�-�ڸ����3��Y'j�0�|����0�+�ĳ��[���Ʉ��|n�9���s;����0k�?[yռ'��0�����\�c)�K���c�H��d��?;�3�FK�rX��to���[J"�btt����,\��:����#q�8�*}�����[͏��y�md軙��qC�J��E H�j���o�`4� �1k7h�Y�:���f�EG@L�/�U�"c��w�{�� �.�$��	/�t
3�����N1�$�mpH��,�)�)i ��	;`E�Hv�4Zً%:���BHK�%��AN��"n^�"�^�+�2�(~
:���=�~���}R)�-|ĵ�}T�E�)L(K\��G��Ʊ5��

��������U#���Y�����i��Uft�����BX�T��\P��15���=_ǝ��Hjf7�� jp��Ϫ��DG�Z�E1e���t-�VZ�"��6�vdǨ��Pgy�/%���3!{K���KѢ���z[�\H��Z���1�n�!v�Z+8i�{T����,]�2��"�{��rX$pu�Y��޷]���O\q���q�l�pB/>v|\��9X�L�h��+�(`�E̮^�	.��l��ol.�JTh����-F'�Ek�� ��7 �\#uo���׿ eA��Ʒ�?C?_�DP�?P�:��/�?�z�tG�&#��i����Z@c�M�mݑ��^/�EgH2(��%������V�R	)̀��9&ʺ�L�xb��5_Z	6�/	a�y�Qͥ����7�!sa7_�j�Y�cL�k=�COr&�O��E������^��m�.�ώ��n�r�   ��춒�����\��UMP~�d�X����N�����鸟�	k���*�I�������_�g��"�@/1��]�q�tR���}( ̱ 6�!�{�2�(kZkG,��@Hss�a������G� ��]�� 磐-�l���ck%��	�C��ϼo����R._];m~��y_Vu����L+?8CM ���ٚ.�ܧ́b����^��F���C.�R]o����)c�I.3q'NF��@LN�J4��_�`��3b��'�
4�t>է�!��Q0:�s�@{(�tС� ����%)����YF�~�+X��p&�>��&�P/�8dD�"α�V�|9�iw{>j(�b$[M�w���Y���f������k̒�ߔ:�/��qpj(����vU�w�B&9�F�ܱ�}�թ���h�c���ت)��U���L��Z!Z��qU~M��Hs�{�OU�T<�m,7&�Mu�{��SR�c]������z��3}_��t��m��ϰ�w�h��5��J/�1���^n��lwb��v?�yU�[���f�͞�|,�d������Z�gB��W��}����.���i;Տ�wG��=��\-��C64�{K�(�B\�p�c���d�4�?eQ��<����ɔu�ц D�
�o�(K,R����km�_`x�a��H}[��g]#�rְv�v`N����×��7ik�s��B=�x��5��^z�@C{bi��ñ8���� �V�F��:�(�Y�����g��6L{gPo�f��nm`P����8#W{t�mUw��=U�<	aݺ��3y�^���ύB�	=�J�'y9����������>����\Y ��
bp�mC��L�����WO/�����+�f�g0_2��l:�@Uh��Ӎ�yDc��^J����6�9�Ѡ99A̠垍�Aj���$�t�\ۦ1�͢�X2�!>ʳ%�cX��}k�TPV�ή�p�4�N	�΃�|�����Q���e�
��"�GՉ|�]5n��b�̗)�S+�)mh.�l��5�g��!S��J�m��Ϙ�X&mT6�_��j�I�A?ȁ2��;,S�f:ї(t��I��7��jV+(���[�Iq�"�G~�z%%M����~ⷮЇ�:l]8��e��&C�j���l���R��EgՓP�֝Nso����MR���7���ӴtXA�~�M(��Q�TT�+2� ڞ����,�a@m[�R'�S�U���&*�;�y�1!��h.Q�z�H��0������o2%�yA��;L������DmY�ipoߛ��7Y���;ɝLC=�*iR3�d?Gn�o�+��Ş�� Q�]hpA�
�̬���V͔S 2�^	����,�}I���:-� H�o@�ܪ��>I�f-?�K ��ƿ? �.cs����J�+14�nģ������7Pk�E��L�ǲZh�0�Yă-���-�r����,�[u�������Hu��@}���)
�!;�D��帷���'낿�:�a�=��u�v�-�^gS�qS�y㭆�[�L��g��M�%�lV�蚪�]6S�-�ޚG�ڭZc��XUkk���]P+>򛰴`�#�,�p��.�rӖ��)Z�n�@-�6C�̨�G%��c&�I��o�����m��5Ш�����oA����i�`U���D�<f�xh�  =s�r��
�o鼒W-GT=��h�Agk�],�9�Nν;�1�6孉XJ�������yK<����ř�l� y�w��O�-�f^>՜���QL�G:SJ]��Y��v��~�hJWr	��ç�'�`-�ƮF��Mٴ�З���n��Mk��ˁ~o��u�:�[J$4�O}�ꫥ�Kѭ��J[�vM���O�F��/� h,�g�[O�8���w�n�$l��G��tQ�'���d�y5�*m���|���*%z���ouJ�qz]�z��s.���EN^�P�<R���h��!�3���c�[4����3CtHaw�O �����.��7�D�ߴC���H����;��2�n�E��:�޴��m��'(��>���"�v�o|��k�9V�~=�����A�;�D?�`.�IK�����zԎ���W��^�z���5�y���3^��W��Z�� ����R1�/��ve��%����"�@��6�nݔ���H�s�*��{ �:znmm�z.h軰�������8�$��h��l�ޘE��gaia7yn<R�V��pF��q����a��q:0H�V,��Q���m����e9����6��~ս�J�� }�	���x�0^���\���_���T��G��>�)�bK�M("�ssR���l��5PYՎ�T��*���ų�6öQ��y�F���h)!�A����
����"�:�J-��4�`��p�w0�e���!:��a�?D�(v����#:7��֮�nj��<�:������[�x"Ҁ�%=a���t�Q��y�s����SR'e?�����&/�ha̮���Y���؍�z���~/.�wt��x��c5��<;����ҚypՁp$�)>%]s[Q�^K��8y�%!��j[��h+ĺi;p�}��A�r��b\>g�=w����iwr�سa�m�X�2�εO�D���$��v)�k��c9.9�z�nL����r 412��7��H�>b]{/�k�g�@��q�(�a���9ƟRxu��s��&��&a�xɻ�`���}���x�y���of.��+�|~!���J�-��Ǿ�Tg�����S����X �:�p�W&G���-_h|�h"a1 �l,��y�+�)܄f桡#{��5ɬ���w���~`�� ���VЃ�v&$�h�N-�ž l�}hf���r^� �k���<�c���ӏ�'�u��'%"uh礉��5��Q=AfE6�H��E��s}�b<ͅ6�X6�"v(�1�
<��Ź$Q\�397{�զO�E�p��i��r�=�:Y^����Q�,�KQ̰X�q�(�b�F��%d��Y�ʢ�7uc�������ϲ	��ē�ѳ�v�Z�!)3m��F��x�lK�L�\S*G�<0Qp�z����X(kq:5@��Ö����gp��%|�9�팥#��]�1k�+�LQG��{e*7�Af�,�:$h����Æ���b[Ţ�O�#\MQ�oV&U.�L&��c�ФfA���i����D�mX�٩�rnMp�ݹ^�h1�M�rփ_��Q�u��$^���oa�DV����mS��	�E�j����vx�[�fR96b훾QW����Z�߰/V;�l�\-�I/�	G.AzaI�\��H`��~[J[n)d[~��C"��X�h��Ѕ/6M�H�n'd[VA%���f�HBo�z�tE�4XSM~��+�y��=�+!���-�3�Pj&�11��]H�.g6�ȇ���ho�B�V�6��m���Qm���Y���1�њ��[&ӱ¶n�v��ȼ��Z�L�J�H6;�Ct?7	�)F�/�.Ժ��f_{���E���˸1f��o��e�*�y�D�F�X�8������DW���}�� uJ���칦�'j�ٴc|���<M�D�_�g������M �������_����}�w��Me%���t��p�����__�
Q�9š��FB}=+c�Q��H��*a��Hٯ�>��Sl�LdJFa'��P_8��(�ʣz3�U<4�@S�M���G
�r;���"�q�nrꩄ��������wJ�l�h���'����J���KtQ��|��=Vw7���H}x/��'��4^"�C�y%��oG4:���+�:�^�؀ȼ�j&p#:���h ��^�9�rM/��:���,��:=���o4:t��_m*.�nڗ�t݉�Y[	�ܐ����B�Kܰb��3�o��#Xx{s�I��0-:^��JW�/ύ0���k��1V�G�X�vRKI�Ka3�@�?��DZMn�_*��D�*�_�t?}c�eȀ�N�'קzנ�n�1Ā9_�)�D�X�o���P.�SL�S�C.�0�kHhd���-��J*��qu�F��H�k�c~��Ո�K�	^���P,�*3�h̔)Dr%~����-۲�]Y���E^�2��E��)r�%��.��t#��*R��h#�ՔVR؟�| ?ɕ�vH�E!5w`�X�M���$Wn���-���&��ø�'�`n���8�"�!��޿U���q��F��5x�o��t���a(v8�gb�I(���ǫ���I3x��^[�(�v�^M�/��d)�b������Y@�&R��epʃ��(�*���,k�@&�i�i�!�2�U��r���T�8Ǘ���p���H��3�f��/%*e[��J�� 쇬��GT���5�n2���+ ��s
e*)4�2��2��gx�w��>�9U�=ׂ��;U褛�HTS�[�\2&I�����T�ebi�eV9��1W�������^Q�d�4���{��*Q���ۏ,'<h���f�~��iJ���إY�c�C`3L�<`ő��Jnʶ3�ɶ���6�Q��C�#fK���	���0T��[R�'\Չ\u��xe	��>�u�Q��n+*�Qb�n��ި�7��4QA������ױ�_!m�T]��\�B}��1%�1�g*3w��g��lu���A�r�${���떍�1ЩR��{O�)_V��Hߊv��Z��n���λ��^zߊ��O<��MW����}���,�O�����a5Y6#�E�f�}T� ���
����ۙ9��Y�^j?*��TQ�`�-}N_��஖���# ���& �=�")�t; ��J�i�m��i�������*�8usK�����FEJ i���D����dP��W08g꒨�����G�β��*����eL{�$#E����v|R�� yBk�a��|� W�;G�z=���ˆ�J�2/O�@=�']A%�u��9(q��PkR@���p��Y�`����lb$�`���+xr��='J�B�k��V�W�U�g&�m]q2B;.׵�c�TT�ק�i
g�;h����e�k�qg���!L=��W��_��]��o���/�Hˋ'��*���"��(�Y�z��s�>�K��8�������p�	�zuO��-P��@�Aw�A%�{ֺ�B���"�߰E��[J���!��\D�6(�$��N1�2���� [-�o@�>�è�o��n���Ey�\�5�@�[��,�WgU=�G<X�\wZ��ɐD��v��#s5�34$����\�~5�4��L����pgU]B#U7�P�m�ߗ�+ƪ�I�{�)��Ō؇���H��!l��1��n�_Nx��g�~���$�/Ţ���i�����e%5��Ik�t��י:s,�L����h��8ɕ��I�B��p��g2��+�q�`6�4��q:��ZJ7��5 ��X���qK^$��M�%@!��~�a��9�Ҙ��++�_�-��[/�zИw2��<)\��Ox	����M,{�F�֪�j��Y��--����{ݘF���!�� ^C	���C��?><y�+��L�4�lh�6�@,��ד��AQ�2r#e���敞��3�3>�үZ�'���
�2Y�2����TQ
m�w?�������p�*���k 7���1�R����\#+y�H��&�'�r�]��S�q��vЙ��N��N�F����W��#3O�ۍ� S9�9i*h���|o�`�)�G�;�g<��{1Y�T^�92*÷�>�{Q�m,��+��,K �(�d��×w�D�J��.��9�6(���n��}i]P�J�;\0�o�T5�8),���_v��e���Ά��O=VG�޸,�P�&�X�c��KB�~�
���r�{�M�/NB����#��/y,-�Rg� ���I_���q���nm,o�K�?P��t_�>`��ڎl@�B�ӮZ��D��Z޷F�p��l���ahÚ����^M�;C�B���l �'�e�0�G�#��-���_��2ԭaLWtղ�	�u�ih9At��VG�nhk�ǣ�-�ν)l��T��t�>R��<�E��Ҕ2�<�$�Kl=�t���6��Ȝ���͗�]濩�N$}*����Z�~,�eSr�<q��QH)�Y��1�V	��ߎ��\^4���:"�Nj�#�D�c\�a(�����.!��$.u�k�t�.Q�|��o~E�J���4�K�J(�枋U�z��-TVs��㒘��B���uI�Q�yg����H
��^����|���}	�{��l�
��Ġס,�����s1�F��0g}N ������������H*�.�P�߯�Bj��t��z'�"��HA���2���w���;`>$F �"D�փa��c'����P
4��<���)/�W|q�]&%?U��d�.mb�.i�.�!5Pdm&S���R�x�S~����&Dsaə���j��~��sC�L^ϔ#����/w%�T�-J�|>��x��k��[R�� �ZX�䩀~���hl$8��A�F�N�I1�;�5��kk��o�Bd����u-�k�g�!xU`d����ݚ��E�j�Lk��]��i����>i+��<�4M��N���\�L��<)c��H�*�p�9�q\��D�6�!���L�;iKh�U�G(��5���پ������ݣ�EJ�1�R� �q��q7{z��S�@)��� �s�&���c��ia���,Jڝo����4�U�nY��JS��f(q�9A��-���w|�9��24�_�V�8%w��#��+���ݔ����A��$��4���m��yd�ɛ�;6
ҏ�b��SQPu��H��~)H< �=<��pS�:�*��-�ѐȸ<$C�m{�BҦ�F���͢i�E�w?t{��^�@(�O�ܹ����
�n+��ڠ�����l@�L�����E��I�2P��C9ѓ�*�wt����}�Ȳ����;��	�w!Iu�_�7��¾V����O�C�:��)����_^�t&D�S�4�(���m�Ǽ�#@�B�	�O�z���r�'L.�<�sʊ�8�Ͳ2[kj׋��e�H��gT��'��;�<��:���N6;�!IEh~�%�\�|촄�a�u�A3�B�Hulv��̭eqf�ל�6��C��i���R��l$�m�׉��C�p��ې7�&H���Х�
����Č�ju2?��(��yE0��2&졀��������T����a*fX�'���c�F��f)�܂�p��e����n����e&{Վ|�?W�*�Z�!R�T��(^o[L[F�I �a��Țt@�Z{���b��ǻzU��!~&�h����eP�w/,�J'E���$�վ�$]����Bړ�2�YzS㚄�����Ht��)�!��������߇-^S
�<P��R��(���EDZif�\�)lTXk�����@^W6 �_4�\����(V88ih�4@�N:��8J߳O�- *����# �6-�ReӇ`D��C��M��F,wܹg^\m ��^vmluC_�? �y�29s����2V�����d�_>ɾX|�#����ն�1�3T��IО��/:������\7hD<J���P�V��UvM�>g��B��C��@&�����Q�)��Q (�bl9��ъ�x�d.��sZpج�E��o�$��%=�_����ʍ�l�狀OS��d�f�p�����V�3�"��e���M���3��,C�8h'��~���Qk�e��%G�U�r�d8�Uc��f6+;E�m)n�����B����&_�G�wH����-���.8
���K'�7�SoG7����``�X��k�|��>! o]��r����S�����al�#���;<�<�����Hw��n� 58�;��ʀy�͵ h����M��EK����jt����V��R�^�;YI��gLJWUc�)S�3�c�c/p��W�P9(��L%����̆/� ���ۨ�]���ITj����Í��X��_�r����Y	�$�����Ed���]J�c���9G�,}"
������A�A��͢��Z8�����F�[>��]��O][H��X�5�Oiڭ�u����F�.Q;����"�d)0��4��#'N�b+��/���8���˧o�"7뭵�cc���P��ts��=3	(��5�զl��CHr!�sJQͯ�0q��[ڎ��hd����Zr&I~1j�rr��)��˧��^=�GI�k�=��v�@)��0��r���M�hه�I����4��X��Lt��gzdŠ�c�;r��Z�Y�P����(
�l����/x��mE�މs��7,-I����d��?YK�QΝ<���A؍�m.�!>	,%�+PqK#��N{xGp�H���H�0�wћ�V^��X�=X��V�4Wzh-`kn��gO]�� �nw)t�]'A%-0�T�d�������/�z5+T���I��ab���{����f���vZ��^��d���M� �-� �$+���3mzoWL'�k%r��ˆ�l�N܀�u*��N�Yɐ>�E��^~�u/����>�tt���ŝ-iC��$����~u�kz���1����"�6����g�z�9j�@͉���?%�&T����A��g��r������P��-sh�
Ʃo�*��ֱ�:��~���	:���V�C+����/r�N��&s�Z�	��q�0TApFE�_�Ώ1V�O{Kj�!)&�:w��315L�R��C�����|�K�_��#?��x�IO(OE�ʈ���YEٷ
����չ��x���.��>s%���%E�;!�����T����Nǟ�D�j��;2�)	)t�s��UmvdV�++�X�l
�H� >*1�q(3G]�cCJ�G�<F{�"�9��Q�g�p�3�7�mQ�(�'��G�`�Օ��wCw;n�5�������2�N�-f��c�v9H�B��`���a�߅�c��RZ顥�=���&���K`����"�>�;[� �lz�xr1�H�"C+��h����cu]�F��@�V�z�0������{nd���癗�LUAp�cD�.8b�/g�44���������������'r3��`�V3E">��tE�ϗ����6Y�0q��JH
~Ėl��Kx$JcN��)�Vq�{��LD�>�@�T��^��=t�s�ᇆ��ѥ����M�:������t�<��N�Œ�[!A��!��?G��J�������zL�|b��M�K�0� �������":�w�#x��VEL��o�U�Qy{79���,w ���@�k����TB��U}�J�N�wz+4P/�e5���E�>��ŷ����P�x �w��P�n�R���ʰ���]��'\L5��d����R�X��;W}������sg�<5˺h#D�ab�D���d+�����d�B��w��@�'ow�!�m6���=��/V����Nd�=
�Q�NA���=E08���	�*9�Û�D�5�!�'��ԫ�����<�^.*&;5���s��h(Y����JQքb�6�4�:��t�E�?8�n��_��~W���*�i0��۫:u���k���l{��hl���"r�F��E��Н�@*(%.�t)��$��A��Jac�t��+�K�S��sm�%�=dD)���U�)J�@�9�G�EJ\!����L6��a�w��.ڑ!;	�O����
U�3�ȓ�sj�@�W��!s�ͣE��4R�D �T<u��E ���g�����i� �>LP3�������"����L������ɇ^��m�E&��\?	JX���l��5�3�/��Nh�6�}h�)��O��O�?���򀴐q���L�)1��� Z|d�WA�X���d�}������fuF8Un��1F(�]F�w]d�������s��G�n>�挹�Eӏ��xAk���yܰ<"����f��ޒ,dF�"��_s%�����p�Z �E���`�2[�P��t���o)Ti�uLk|-Q��Y�U�#-��qP֚�9��Z�۫��V����ek�CB+�'M�~�DI�$����x���{̵��a\�>�]G{���|�XQ�u��?lA	y����t��9�n9��	������A�������[�X+o�ͨ߃�U|�%��d*ƷÈ�Y�����J�8o�ՐvoU�������+:d�@���JV�R_=�R`"u ov047�o�@L[�
��7(/'�ݫ�R�,��_`�C��)���&�	�9������&;O8�=������pZ�+O�@o[̮��H�TP���F@=��K�%LyW=@O�Vq�=$�C�(����^y0+�l��͞8�3'�-�-w�MQ<s�x$�CZ�Z�r�(2�'NG붬X_mx_�0U�R���D/w(�B��{�1f�J���Wߨ������B����;%x<�U5�*�5%w��$'�Q[De�Ӧp�P>5I��s�̌1D�xSx�K7�^?�����q�6b$MAr��/��_�*>�#޽��f��zOU6qT�n���gے�K���)*�m��!�ҭ%�,=���=��}^,jm��:d���2ؕ�(��$�̉��B�k�ZՅ5�L��s;ɵ`k?������{��@���K�b�ώ��׻���	1d�),P��{�h�a:�.i�̩��eG��Y�&��hWR��\���m�6�*  Iѯ@[�r ��R� .~���fԄe���1P�@�j��?�U���F���(���&��N��k�r@�?;N��4I�5UJ�[�t�؟�s��J�hk�@�$�8�sL:lkC~�W%د�t���,M�Gա3zT+9[�u;",�ظz1S�vV%��l��߯����٫���d2oK4�,�R�K;�*����ݣ�dV��˲�z,3��f_�;ԇ^��ܞ|��[��@'|�$�����2ߨtuEk0�I���_�-jF6�Bn���aб� ���3� ?o�x�7Wn{(^�jl���7���"��Y B4I$7�d�o5k��k�$�6�<�O��&�}K�c��-�?��y��	ӣ��fϳx�t�hk���c�ź�XC�ڥ�
�lD}�D%�C,�?��Q��F�Bi���ts ���1��v�0�PZ��1Js�9	�V�=���"bw�(7v�4�/|<;q*�$�Q����i��
�s��b�<�Ğ���u�;��Q��"�'��q�+GwBD6���" ����,�,}%Y�XT-�������0�.����a�Iu93C����d��Rf�H,�o��E͚8@��	 �$�lU��G��=��`UwM��C^ß,���B�ɡ*���1WIK�`̉e)�Ca@�2�/���"��fd	B���[�.m J���oI�Q� AK�i���׆f�s���������Հ��P�p܁���͌����|
�ķ��P͔�S�QQ�r6"�qv��E�Y��E�Xc���tĐ��yζ1�B\���r���}mP����V�c�C�q��YZ�by`�Z��Cۼ�nxa-:tڳK�����vYhw���F�����:#^�Ӗ��}#$�l�0 �A�=\�5"�lù��ƥ��n�畇Y���܅cg��T�@���0F��M�J���H|rD��(�ve��ġ�>�qe�,����ܖ���M��v��B��#�V�\�7%�$\����b��df5t�=��;+�
$R���l���9�����n40G���ӟ�?��ъ��Jp�v�!*�ՙ�q� v���sBU�ӹ�4�#7F�GAf����V!�Gt0��Ӟ��(�j�	�����H��_뚌� �&�zh�����,�V��'k���������$��|�Ԍ]*صTNr��mp�Γ�����]�Q{v�����)y����Q�����
�>u����~�ɖK!��Ӎ"o���Eә��T��&SY ?UˎF�b�hB�wV������$:���N�|�>�F3�ʾ�d��fڬ�_��ؽFi�8��ϢUK��W�K�/��3�s}��U&O�آ'��IT��1�1ć�pr&a��n�Ɨ�8,�d�%��3l�`y�p���k�ћ�Y6pFg��Uq��ٻ�MZJ[��/9�56��u	C���D�g�Q���S��ڐ�A]q���×⢇+�r��T\Ue H�<#�7��oVH��({���	�/�5��FL�fgz��n���Nf� �5��Q�*o64e7{��e�����}�>i���;Mf�.̑�B��9_Ԋ��5Rtfc�\��|Fv��5��_�I�'�Q�ĺK/������4C_D�E�e�<-���k�}��G蔫l���ͯ�*q�P���V��<?�U��H�+zW�W���\y\&�%��=���j�k �d�_��h=ˏ��u~�怦���f�ך��1Y�շ�=��{�C$p������>e�XBCHϷ�3~KkT�g����k@��(�{כ�/ɺف#g\�m�V����[�EPYL��5���)-�8�f���\n���f����A�!7&Aa-�  U�T[����w������%�q=��t&fۦ]��g����e�1�Kl�֋x ���+RMz��.c����xF*�����ۀ76G���#�Y@Wt�H��)$���R�ak�X�R���y��E��`�������o�����jg�T�Gd�,����#�0�Y/�0�$uX�\�=���ίN�8u�\Y�4����P�����t��āq*��X��̐�{��[����گh}�c��Ѕ��j4P�!�J`N�M�ʤX�p�IZ�:Z'3D�/����%�+�_�@�=��& H��R��:K�m߀L���R��8�~^I�L�jm��A�t��WY���܌��Z,β>c�NT7;�ljWHfڻ�9'ҿ���鯿#��R�R��l����}{��Y+�cxf<�h�13j4̕�W؎v��'�! ��v~z��H�Y�-_�s�#nY2�A�A�}�ȑ
����Yv��!��|O��o��15���֯�e��~o"�6^}�JL���81��-~�������%q���j]6r�4�׿��[�h�F��ߺ>�9I�/��JtR�+K
@����N���p,�o�!8�	(�z���gd����S�(
�|H�;�fɩt�z�������:^� ���p9��t���7}���%���OS<xh���:uv&��u6U[���޿J����x�����DQF�����V��t��I�SFW�_l�.��R�����QQ�� k���{8B��C�_��t )[��5[`u&�u0��^�X�lPځ*�.~ƅh��w�9�j�T�b�xHX�r�ώʯ�f0��8�@�5��:r&u)ݞ��R{`�(N%�~ݑ���U2���� 0|���w��}Α0��[6�t��1ff���+���	
��2��uI��MT�9���4H�V;9n�&�Eṕ��\��kk@
�]�QI�;u���~1�K-�w]�.�/�3ޛ�XMR����Rf��9v�d^o�  �'���?�/Rz��<�s������퓩K]1?^���)��~9	��?"W�ds:犾�"CkcZl|%�W�����'Fl�f����j��}L~�H��3,yן,i�*��*�A˖��r��lv ���^����ꏏ�ޕ�7�CR��k�����M�8�*,��a4|�d�/���� U�
����:�Y���aK�����鋹�Ē�t���LԵS/�@�����[�����t����g=]�������:"���/n����U���y3�a���^G�����]�����/�I�/��"�En���7� :u�,(�����X\&�t����%3/c����;!-��0dn�/-\������_��\��i�@�/=},��9��J�N�cBE��*3KjbD�x��HSz�]�#��١ɸ�9�'va�R�Yi]�?�5Ñ�r�@y �n5-H�J�ݛ�ڷ̲I|S��%���M4|h�G����gr�"����:$bb�R�γ����J��G�=���Jq�����
i��{G���P�l�a��|��jy�J>C�p_cI� b�I3")V%y;�ґ&� *u[<����^�*�Wg��
BOJ�Kr��:�%E��K=
�:VFa殾$�h�ùz|������u�}���Ϩ�LJ��ѵb��8����PLϺ�)t�$��t�E�0���f�<��Z<m�R��+��-��"�рm�v���e@&NK��*x@ĸ�Oӧ>�,��L ��0�@.Q&�p8����PU��REd?��O����"�TLW����o2��m�(m���wo�-w�D�%Uʆ��n#K�_���6R�!%���WD����p5�>%�\����)���}�~=?�Y�ڇ�s5=�Tp���������g��<�@����ʉ�O�=Nj�Z�$l�w�D�J����B�?³mK�-&L��;�� �s����t�u���]w����V���� 3n��Z10#zF��R�̇�U5.�Jg7��"�.��Ɵ�ޓ����<@������N+��6��{��5� C<��K�yr8�|]Ņ��5��N�{>\9���&�S�X�O���B^ �̧́�ۢVe*�nE��m&��E��^]�Qg�p"M�Q��QYGّ�xi���w"�8��a�
/�/��R$q[ 3���ݤ�@j��~O�6�g��S�Ô{=>��؂������~t�UZ�����O��S���sK�Z��'������`;�R$|�O�4��������OU�ϩ����a��.�5�ZE��oE�� !c�0��U�NQ�u.m$W/P��� ����bg���I���U!��e�o�%�W���������(�~
Wi��_��.N5X�ب_1�qb�M���ȁ�+⡿-i��{�� ���E5QC,�}>-�3�-u&�,�U��2+�&՞P��ŏ�oZSE�,�r�� �D��u/�exݙ�8�:�͹��Q	�|��9�
�|i����/������B�c�v\�Ȟ�FZa�3$!�&�S�� 1]иs��*��WsN8 GО�+3�
{�l�B��`2���<;��y��m	�O���Knm�u1ukK'�z�`�[��a�	u�uh�Wt�܈��;��5dKdR�DC`&�Q���x�߆�R;��ع>�ɕ.II�.g��*���Ż�� ��qu�&�Z��g�=\�I�bç��Ma˖�B2����Mx�A;7��O��0df���E/�"p�3z���c��Z퓚/<G�F��>w��Re���	l�Z!P@4������l#릅�1ޑ<l�}��U��ke58��8ؕ�~�=��V[W��Ӓ� ��gD���ܳ��?Q)d{Z�O�r�K�oxJr�	iqd��T���D���caV{J�G]���$Ս�Od�Dk��֘v:b��4���M�7�$CyXO��BLN@U�"����d�9,�[�yE8�2�]C23�F?�@' c�Ug�&g���^�S!��,�w�IDC@��t�N3fúQ��� �r�����=��<��P�����n$a����\A	v;��g�D5�R��1�5/�)(N�Y����-a��\��#GSĬ�$�]���Љ<1�_8<ֻ_��,�w�`�W�^O�A�3YX�;5�kq�F�f�Y��B<4�B��j%l=8{,u*�J���
�U�?%E���P06������j/@%�<�� &����F僚9F�D�����Z��LS�e����ޗ�zJ�_)�n鹓v-�(�E���LN�CR���#=��FN��N���-�@U>7[2,^.]P���~|Ϩ-+�{�^~r�Z��-���߬/ʄc����������O ĕ�bPV>���Wh�~�M�� o�f����}[�Q!�����wG�"&�lu� �Q��4�p�����G{�$LI�����z>uL)?G�����;��r�9$-��5~��{|��e�aӜ�	��������KD,�*��w(K����Nǔ�o�B@�3^��m�D'�u�JY����QC����5��#l�{5����6�?���abq�)*�P8�}�lK�&컣�"k�Z�r>��d���S�Ӌ�l�y��~Ah6%�O�v���mѳm�߀� )��X%g���K�7ʛnf.]luM7M���q���k�N6͗���'P5_�)dV+f����b}�&I�����"��L�p��*I'^
jl�&�6#Z
���j��UBUS�� N����Y�nX��,hC�z�\�_qE����>A�;<����!�t�\MPC���92�s�"�@����+�`��w�����%��n-�J{plֻ�~�QH���#|�G�R�QU��c��.���p�H[.��3�$,�s�u���S��\���6Nٜ"^��I5L�P��)Q9�GX������|�q�V�[rx�l��$��e�$گ,D!��3;��_�.H�K�([pq�[i^�,��������@	u���w
^<��ʛg��so|0����P��g=�&~��Q³���f|lWF)+�8՝�<��K��!������c�G����[�%�#E���%"��v w�m`8��d��>�dT�1�zAn������j���pCĻ�H��Y�h~���&�����(G��[��h�p���B��A���[�]z\D}ۀ��$j��t��]����<C`6����QP�`����D�:���V��YV{yΠ�����j�8����q3�V��u4.�v)���q�8��=�K��>�t�4���
g��ń��M޸O�)��E��O_m�@� ���h2���:��A�-��l1�,��E�o��zפ ���>ld�����Ax31�K±\�����U��p��mGD"���ڳ?�(��p��0�Z���*F]pxoQ����� ��Y?�W��y:�z�Q�i�bu��Pb�
�95�}�<����:������Z5N��NBSx?��\��d�O$97���4�ǉ:����@.��{::�<����I?�C� �"���t0KHfɵ��r���.�BK%Gy{��(Z��(��QR4W3����4rz�>���m|q�i�&pye�]F̈́�s(/�����5W��D=�?�Ŭ�K�{��7�F,��4u�Q"�����VbVTZ�2
��QP�%bg.���vZ�̓y�. ��{$�xK!KR#���r�4���%�d����D��n������TcT�������=i=���`��X�~�����ؔ��B{@�a�[d@T^��;U�2��mWܤ��*�u4�z���8�gF
?ɅP�%Xĭ�]C\�^QX>?��)��I@�2e�DfE/ɩ��m�(�=�r��f�m=�-��~�T&�^�)��뻣��Ĝ ���D'�r�C�h,6h�DH |ӆ�>����y���oU.���Լ�:�US�,�r�&�gц6pe���xMQ�@��Ҹ������ۆ$�m�z��f�[�fY�?��������ۆd��-�|z��,��I���W�ѡ�������d
��
��R>&t)�q��VXR�!�ĕݫE���o>������:;gg�֞D5m'�I&�&�Sd�4����{o1�l�c��wp9��	�����ƕ�����~fnM/\EZ�����s���-h��xk�9��0�%hZ�>v?%��u�?R�)x��AH�^��ٗh{	��uqS�I���j�T䯙t���V(^7�W���9�>�;�����s)5T���� �s�)�E�s�AsMrٕ�:},!b;��n���e�dn�6��Zl�C�*�k����|�ԟ'(¨�=�$�}��/���q�1��-,}�U��f��r�:Ҋ+ T�N7��|d��y͓+���7-:���2`|w��������A6�̉��"����'aPg�-�趲�:�+�XeQ[U�{�\Nt�`���a�s ���#����(�PHiÙ|CCN�\l-��>qd~�, ���gm��3�d�n�=���],��F�>l�&!��L��F���wp0�"�P�9�]:� m�6>�`��-�C�2��l�$g&R��`�vS����G��2�n���{�%QbV��Q�10W��m�SU�t����m9��֑�C��,�����t#�Hbg �#������@
��.�v��V�vbt0R{T�ׁ��5TL�a�0��!��ţ�ߘ��CKPo�	���5.$��i�6�.[<_&��N͌�&9<8��܌D�I�|j1v�eݰ�G:��IA�Z>�����	�l�~Q��!%⇈�Z�3	�<�@+('N �̧|5â;N��`��J��&�N̨�W�s��Dd�	3��3����)�7	B
'��9�ܹҥ������\��/��0��y�ɜ��%
��H-���� O�!�N�UY��T�k|��P]V���0��0�@RCv�8��w��bH�Z�!�#��1�: �v.x�	2Ffj̹�(�q�\w���GS�<Q������� v���u����Ř-�-m��-���B�F�����7��#�f�}�ԟ�#�v �!}/���_�'�6�.�MH]Å�"�Kd���@�i0S.V����t��&\Y!��{_	Sz��	�s��Q �������g�4B,�� ��G �t�ۣ:n��s��ŵ�]^���+B�dh��������ݽ��E�u`��� ޤ��UT	��@!E4��~~���]_9��+��p����'�(�/A�5���|���:���X�݃�Y�	G�<�����I~��.�n
w�+�Xs����Q��-<^�7�hS?���yCK�����h֛ ��S�'{U��P[�2M$)�l��M�*	�`Ew�x��uRr��G}}k�p�W��ަor�~dZdnq��n�箱��_ީ�&?fG�<3�4P�������S�����՟~��Y�fk
������?��%.b�Ɵ^��
�A�B�{��ok�|tc9P�^���!�Jo����T��|p@�L�S|�N~78�Jym�|��Z�s���]͌�w�!Z�K{�ylܐC,
�_e$3�uA�I�@�a���*'�RR�*MXyLaY���.5��k�[$�� �]S=a�ۏ}ki�LX�>' �Z�$�"��+�;ۡ���Wv"J���W8�{�UUW���
�)M`J�,;��*�{�������yLl)(��}��͎�N�?r#���{ʅ?y�k�}�0{���'#�5%���51$�ضP!X.;T���4�<�����2G�w�಄�D��܍���QfQ��U�J�=H��|V7���Y�m+���\�p�0
���.�w4uW���]l$��O��f���W>�H͛�>�=ϛ����yU����7�(]l����|�# �7��n$����'�kl�l,4�)R���7���W"u، ��}*�[��ǜoMgkw�S1``��^�qQ	-��[�{ı>����F�u_(}miKוT����d�(@W��7�U�h�B�*-6ߺ���k�)ͩ�y�A�[pu�u�'hG��V�n�usg�d_��p�o�O�h�p������z�fWF�]��>�����
hYdTe�ۇ�����[����.?��+^��m�'�k#
��K�7�ѯzF�u0	Q���D(Y�����v�1ř_u#�:u��� �2
1��I�doh.�යT��75J\��b.ɇ��¹���ւ�"�z�;Hr�jέ#�+t� ��?b��1��G�Y>$rk?ŭ)�6a1�r�A��a	�������)�%d�٘���'�����ؖˁ���_�K�ϩj����`�5�zu�	�䁘�F�!�>�)��#P��5�a��c%\���bxx%�~@r�Јf�(3rQ=�&#�Ŋ�d��Wb:�H�@�/zX��]'3���e+����*Tq[���s�
��(|R#�����[����J)qy>�I��[R	��琗��Mܛ��<N8|�~�8������6�T)@�U��Z�����{�9l�>�>�ν�f�"FkCJ��Kr��	8tNn��n��>?'�����ID�Uʋ,|�o���M��u�|.��S
hc+��X/U��lG8�+�2c&�Z:9�ܧ�	Jx0w���k옢ա��$������wx�w�u����J��؍�ˌxQ��y��9)�m���7�����ȹ~H��V1�֮N�Ƭ\@J�,!�^���P���eN/a64޵�����O��\�5�Q��>*p�����o�4��M�
��)�)�5�K#�u�ٰ���-	���&.Z+Z��M#nM��u��7�kAh�׵����3��A��j�=��	�6Ȅ�M�c�ki��v/�xf�ύ���7�=4��!�Pf%��9ۧ�?Wv���;��T���_(�W�:��B�h�[H~I����Yj��7%r5d,qE��r��Q��9_Gg2Y����W�o.���]ƹ������T���zYGb��J��O")]�h ����lv��p-���l8:C�r�ڃ��� �$w�ySƑ�L ��oG�&���hm�#�~�k�`��,����x
�:O*o��E	���M�ZVHd^��VT�ײ��)��cϱ��&���h����Pm���MW�L��̂uAm�ē�_z"̽��=��wa)H:�׹(��',�m�w�@kN�����)��G(��~�+o�I�'v��Y�F�ħ���MJڦ�c�"RPy?��˭u7����fa�~��@p�ҷ.��˷����ߥ�b�D���o��G��3�s��	x�+��>x)A�to!�/"7�� A��έPgM���s������Q^���+^g�G��&n��r(7(a���ǣǥ׏o�����Ț�
���p�5U4r(a�F���)�u_c�d�0��Jd��ۯ�z���*AiX6�zRй}0�|�
�3�AoNj�c�Ĩ����iǏX�����7Xŗ�:q�,�`v��K���Ȋ���ޘ��)�^�`�d��1`w��짭���(�s)�۸T�^S����Lߪ����O��!J�c��䱷m����a����M*�2lX�/���}OM�%&���J�q�e���q\b���f�|P�4|}E@@�	�{�X<Q�L3�K���ǃ�b�ctN��[q�N�����"���4T��o4[�m�3�C�L��o�	��e~�\N^����Z�A;D=ACV�g��u��M�xX��"��G�2`,d?����n����T	� `�	�e��nҹ�R�����_��������?�2�T&O0�D�5XRT3����j(��~���T$�f�rۛ��Kҷu�i�7�`�����(�6��h�V��d`�҇���{��r�Ƈ�6GF��$��>uw<J�U���L�K��|�8aӽ���Q1}pg�^����~ӟQ�J��X���6n�S@�A���E�mΏ��&�!���;���6l�n`�Y>T94|�Rt ���-0�1�g�'qd>%kq�3�F���?�)z���b
�y�(4%]�w�Z� ��;N.2���M�&����<�泼�	3�|��x���an�K��Kg�߸�ɠ���l��'G��aX��� ��- �e=Zu����Viu�T��A$~L^�:6_[�\�F�?�,;AI�t�6��۔��������n�T{6����dD�jޜ����Xi��1v�kx��[��z���鏍�2`��'��ChHvˆa�f�P,�����Զ0J��Q���g��72�EG�9�jSņ�b�id�y�p�BW���O3�y[��W��@�DИUI��N�l�>��o�E�L_�c���$zrc�}�u#���'�����,k�*�H�w�+C���J�1�uT��0B�9f'/�\Z�G���5"��9-nw��1P1ƞ��ؘ��N=@��m�X�\3"4=�&i�s��^�n(m,تΚb颍��v�f���)o�'4x\��i(�bWM��d�ow5$�P$�sv�D̍/��5�'y�=`�F_��Go���{�R�S��H~��mt��lʚ\GX���������u����*�������zX��ڹ�7�#/T���2�Ӣ�q�U;������h�k��S	�����{��vs!A��^UCX��S<��o6�z�]���,����.��X3u��h���H����x�CU"�w��\.��)��{��@R��if����@$��6���A��.)[�ܥd�o��,����v"%��=�͠�66� �}�1z��U�j�}TBfU�0X2�<󟽗�E��C�'ʌ.����+�b�m�JϹl]��h��\��0]}'��u_�p2'S��2����!J�34����'v�)/Ʒߓ}��_3�;�i�1瀝Ɋ|���h�8�5����㡲:�����4�^r���!����P,��i��d�܈+��-ե�M�!�����D�`�y	���.�]B�[x�"����DX�L��A7�f����\:��RW�+퀱$oAʞ��Q����uV��T�4a�w��b�f��[���$����=P�zcT��]*pk�@˚P��gnv ���X�6D)����h���s-�j
��T+�v��(yᄈZ ���{ }�&K�˵�?)��=�E?ཪb%�4waK��������J�u1�2��"_���님����������MHB�.t����~�ɤ�Gl�G��s̽Ŗ�@D����0Z.��bi�P`_c��*EeD۲c(w������2��<NE����~��S��^�h�qf&r�����К���"I,	���ü%B��������" �3ex�^`*��o�F|��NyP=�9�=6%��m����T =�|��W���>�sߓȬ^ig�'�#$8\�{Kd��G��.0�X�:";R�_�t�pz����:���4a�]T��B{�ٜ7>̈́��i��
�I�!v�;v~��7�`;�M'�E���&�8Jφ`&	w�K�9��%iI�	��Z�i�������o~���<�ԩ� �8="��oʺ��<�
KJ��Sn�q���V�?^��p>�Wl 1S[�3�٠*kTZY��9ZkK�&2���ب�8��Ȩm�ۮ��3a9D�k	~��Xfw��,�p��.�6(�>&ު}`������}�cW�e⪷K\fv���2��;e��
�n�s�����l���vz!����@3C���t��͂�[�w<����?�6�!T��Ǽw�ԁ�ƴ���Ɵ���8\( ƞs�2h����l{$�(�#�HF��s���-�=�F�n����~'�a�V��)���Fr2Z~3<��8����k�׊坝�� �ѭ�	2�CөI�ǒ��ˈ�\9�!%�t�[d~i�v���mn�t.Oz��s�9*�={ܱ3o���mN XX��L��ba�+� �N����Z�RV;h��ۅ~M �~���@�q�2�x�l�2LW��� �A'��IF���LM"�埞X����Ol.G�G*����c(r&�F�n���]��Uě�f���݅��.�c�#��3î{}�r�Gr@E+'�fw��Xq�~_{���F�B�m��I�b�jF�%��N=�1��}��h��V��񍟪�IX$�޽oD�f"@ ��W����Ur*A��}�(e$$#zY�U5���'�b�@����);��9L�y�05��Rhk8�Sv+�d� �v%8Np!�0O�O��v]d����Y�p�B��ǚoо�=����[�`3���r~���x�v��ό�]���e��P���a���5����f�yoMf}*6�6;�c���v����Q��b��2Q�r�E�;�����|[Q2TI?$��Z9���(��)tcf����	�Y,P~�3��h��K<�4-�H��OQY�|tv�5F����B� ����k$GD��0G9 ��w���G���*�D�%�Y:OD�e�2��_�fȨ�P�m�����~��M���V�g�}���@�o	|dp�n���G����A�Q:0�Vp.);����1��_�8�sX�{Dv����qg"jQ�����Y��T1�h�IO�=�Q�.as�@ir���*�≛���_�V�p��>�!E����$�Q��87 t� ΢�
��h�fZ�W���UG.Z t6�8#�����?�~���b��Ƿe,��%�X��\�����N�h&�e
'rme�RY��-l���QK�Ǒ����0�8*	���;�;��� ��e�e���G��89�)�KT������2C~�?�gcы.\��4ތ�+�4�r"�5�)��T����E� T��7N-���VK�&F�0h�A�`�� ��<�j�w6,�yz{�!¢����,֕�?���K\)�U{IK�p�{�����3�<��~�΅��W� �-�f���$#�8o��0v�z[�#�eQ����P�����{(�9�Q~F�8H;.P��?.<�xX�s��f�� :��l=���$,!���O�@�^�/R03~���zjX�_%�� -b�"�p�d�o��r�@厒C��-�e G'@�'�0%NNr};��ȷo�hw@�د�������� ctt�9�!���F��s a$���k�w� �X�"E�@ZFT�~" \S��^����ݐ�!�bbq�}	��9����w�B��9�����~V�A6'Q"�>�8�}�jV��M�m��/�쉫���?���x:�	F���Uj�)�W���ҵ�,���d*`_��"P��"Sh+^IHy-'s���s]���q:�,�]�����Cn��6�a B����٬������i��P���c���V��i�6Zt�Ű��ѳ�?�?�U*)�L��[�A�we�TQ����#\�>�'�)�R�)i0�LY�	MB��<���')�p���襘�I�S?p���Ԥd���'��?��LVqϧ����KΤ�����O���M(Ϻ1�����w�W'��6VL���;֚y:�	���:���C\�H��C|����`4/��=Q��.����E�մ8y�cG��uV�!ϝ�0I�]e�Z������M���Z��|3,�<+/���I�2�*�҄ر��:��?��ح���ٝ����w,imJ=j6{��	N+��)��ɵ�g&�6��5C�U1��D�~8
2선Ϭ�p_�#��Ձ�S�ʱ��̺aЁ��vk��6.�މ�d��Q�D������Uoc�ނr��!�U�S����ȼg����ol��]�V�lH"b��O2p	�8O=UBl��ȇ� >�^���X���.��K1O�Gs3�u2F��d���G�^Ӻ��HK�0��7�Mjo���b� -�~Ȥ�U��X��0��� b���o9��lP�60�G�[�����l_0�����[�d�2���o�5_���u���#��ն�qA��z!�M�LL�%�� h-R��@֦�q/W���:r,�4N����ir�d�y���/>Wr��~����@kDtX��$�d���[ߒ_��,��W
�pϠ�j��8�x��Ub���ΥB�g�k_�i��a�\�����+zŪhV~P��D涴�sŕ��N��BSM����_� 8oS-�͖���R�$Gh*�I7�;�6�jV���}�@���tN����i��Aŏwě�,>�J���g�2|�]�\e�<�m��a���1�ڑe�rV��1DgH剖�*R�W+��Y�6Ob��Z�hN�L{��l�&߳;k�Ȇ����JQ��L����N��7��Zy�L2�Q�Q�#P�$5�4e?ae��FZ�n�N��83^�'c0�ٲ��5.��b2nB��g�(?+�^�'j�>���(�t��T�}MA��lK"�6���ޕ�"^��Or.�w76��Z�������yS�����ve`hzXK�`*؇�j�0��8�|Z�D6���.C�M�I����XE����zE���yց�a��V�3mV:N��i:̕�ymbu�J �|<��z�[O��`Q�'�+G��ՎhݪVDA��f�h��m4\"s��z�S���`\o�0`�P[m�'��aB$��U&7	H[ݕ K�����	�S]n	�id���)�%�U��-,�^�A�r�+���;ff�	z�E��G�Ҳ9v9���%h���b]+�&dk��S}�Q> 1�T���nh��e�b`�l�
�s�++(�0�[K_Mx�|���R�wvY�xG��� ��SM���R���NeO����h���pQm�,j ǂ�<w�F<���քpķ�!+4A��|<p�g�uw�@9�KdЍ�y��������G�vV�;^p�u	40<�#��*�t�:�^����HN�h�\L�f=@\B��"e��Wh�+�/w^4��q4���y&Q02��a'*�;�{b����2/�4��o�ۆQ�7��/���G\��*b!WM�����#���phQt����k��(w�i칣:�#C	�G�>b%����*"_�aS{�]=�dt��P�}vg	�W�#a0��{�6]���]�&b��ʘ��|���F�5��j9b ��e��'�AT����2�5�&�����<��OP;��c�A0���>�$n�Vn�p�*�G���p��S�uJQ�{��@h�X_�dw3�y
�-�%���L�編��3ˇu$Ix	��^��	��s�F��'���ٵ���S�!tF��6�=�X(:��#�R^��i����ĖL_�o%"��3��@�J��� �_��Q'
���\�!��=��r��;l��U��_.�uz��ZX�+��R�gt��J�����7������B96a����;���>:]�-h\lG����� �%�]�m7�֖��;�D�/�K���WYfC/�.$տ;��q�r�B��]}�2��r�抣���(TggM���m9�σ���>0��R�*o��h���f_K*�x�5�����9�H���(�z�=+�Sݣ,��b~�ϥ�_�\F��-��+h�S�+�Q;�_ak>�5)ֶҬ�\ˋ�"�޷�{���R_㑭�Q�{����:6X���na���LU���T�W��'b�?T�V����s�Gn�E����b5	�c����$nN����g��Q�x�������S��|���o��5�ū�%>ψ���\�%7x��?\M����E�"e�"?=����nD.��*<b"�x��sȡX\I�����5 ��F�X��:�o�iՔg��;5LV���!�!��*�A���F��a�V�7��|i�'I�h�\7�7}A��5��I���f�����T�k#i��%���MI�'��6�P�[��c#u��ċ�%�Q'*T�%�!bP�1�uM�{����ok�~ΏZ��"�[2�i��j-jӐ�9m���uV)�H�� U�e&��rdHWA����?-�uUx�`�T�G�M��
5$����x��'�/��c~���	��>A9����3e�;r���Q�J#$�]WM*h���(��B ����5�Ke�u��tR1���_7�^j\�Y�e0n���QՄb}81��Ǡ�5Zk��E�X٢����y#+�4��(��?>�Ϙ��F�e��F[�'���.��=����ہ�G~�CO�֤�Q��?��Y��wle'A�B�Rs��i��E�l�E���?����:p�ũ�U�U�����K]s��Bѕi�*a��6��4J�(���m�jz���2%�jx�ߢی~�!(8��p>��7
L�:^3-��������m0/��Qtdz0`A�.2��/�s����(ç]��	�����a�d�n��q������0� A?K�U2X<|��=�,#�#z�S��qCГ�?+� Gg�w>R��Y�d�����7�u�q?��ng�1���:�(���I>/O��������l��jhBk�^oQ �~��ћCR�2>Un3l�����^#U�]���$��9��q�g�������ݙأ�����'��n��q7�f��2WN�n4N�\Q��(+2
;��$�B  �DM�L:�b��چM/ѨAHՙ��j��,�d|@#p
�A\�E9@.ML��(��3[0}2�ai�A���&�S��tR$��1��q��ؚ�}X�e�Cdxƞ0n�2�w�C]�oݹ���)�֠T�.gd���!B�d%#�Y��3q񟷶������2���ouŌ�Ƣ��,V�Z]��J���?v��W�gt ��($��`{�{-��wB+u�!Z��'_����u0Q���|�@��:ܩ02�;= &�.-�5Ծ�A �α���m�@�:�0,U�)mŜ�A����N�w�55��ї�S�M�Br5�x=ýA�����'� �to�]8�����8ߛ���2�n��r���+�1^��3�O]0�E���L���֒���!
%�\C��ce��АC>9�XH��Sʗ����D����G��Z'*��b<k}ߣj3B�H���Nab0#m(�x���||E��^���B��Z/b�U�p���B�z7�û)7=~�.�G�<}�6�iX8�e�'�� ��G�kє@^&&����Y	�dȬ��/H!��^��$R���<�\R[�L���3��6�y��R��4=�SE�����@�-w1u`����Ɯ��ɞ�s@oU�C��EX�`ﱓm�W�0�I��Ｙ�����7ȝqKM�\<�w�-�wV��0�m��t������E����W�d�}��X_��<a#��D��f��(��^����{1��$^'��B#���XՎ<3o��?T�����O��qw+U����I$��Gd�@3�����"���Jv��`���Kq��7eS���K.�7����m�g�oA�7�V+ap�T��C�Hs��z{_�d����W"�}�V� ��Cd5�,%��p���I��x��^l�d�yI����lxN�z���k+>>��` ��!��O'���躣�c�� �%f�/�6̋߿�1H��O��f�}̐���D�Y��Y�	O�e�UG�;��"KW���/�Z,�'��r�+M*��A�����D%�F�����������EVoz�8,%Q��'mW�/���W�ĉl����WpE{��U�J)n��*(���߾���l�*|�^eP�䊱hc�m���AW{Q�6� ��@df]2&�f�$�����u�Ѩ�F�5 -;��"�~����<��"���*�q��L�������H(���Y Zx���a�k��K`��HH�)Pmj��Ja�!y��a~���o��,��&�F,̹|�Q����ڽ�����)w��&꒻�'�O����H�������6�`�8�u+D=�����MrI�)no��t���c�E�P-�c�<k��w�-A��;�3�E�惗؜�E������oA�B�|�EL�c%�Ջ
�
�v��� �mz�Hc��
ՙǭ�̔H�6�{N�NM#��� J,��s��fԅ���ڜH̼o�ｵ��/0��8���$�:�j��\���B���up�t�t_�����ڊr�3l����8�ot�K���Ċ�PL�AC?�Sl���w_{��l�,�PS��C�oM�u>����"�������}Ie�A^��	@��Iv:�{ZQ�jlUe�o�zť���;�$RȈ#����ξ�o7I�h:���R9a[�q -J��1�Fi�;�:��X���*^- ��Â�ig'2�XхI�tb�߷��˴y�j�h�	~ADI�F=�/��������}P�k�*���R�{�|S[����)���!5�Q?�HA���l�MeڶO%b���>ϖ��r��|��l�m����<�'5.k?�:�wM��5K�MK���B�k��!N����
LŤ̷}�zR ��0��'��^fp���1Gl����"�������n�U(�㢸Ha�)������ߖ֢D��wNta�b��R&k�O"B�ŲѮ��}��3׾IynT���o��C�%�Lh��N�W�H�"���0�����;��ȕ��~"�߃��U�"c؄4��ys�8�5�ݲ��4��Z�.�V�n l�*VGkX�P�Ĝ;4L��g�l�ҰO����F�<ǡ3��KL�FOP�H����a9�e�����4r߭=������u^M����z����"����6߈����̞�ʒ 㔩8�?2MF�=�߸a��Gԋ��pe���b?��ג�1�EE`�y]�W� e��]�`sԀ��F�����Z��08���k-qw+��~�Ȋ=Um&��^�{2�l^��8���|�p����)�%�+6���qX	�7)!�S�[|�#TАx�lx��Y˔oN�,�m���8蘌���8�t�n��qW��~	�s'eͼ�v�C�!�6��m���1Y�t�����#�"�6���VY�K2O��s4�=e>��;%�CK����u�w� r��8yh���?D8�f�\c�?��p��>#J�Ȳ x�*ů��Lb��9b.����#��:�z��� 9��'k>���\�;Yy#�����FlE�;����pq�gi_Me���C �򖠠i$�rD\{`����(Y�N	2���Ҿ�[D2� �� :�C�b:]AJ�tX��b���T��;�V.��m�Y/��k������J@4$v�^Y.��W�S����F�c��`"���)M]H;����ay�m���q�5hĿ�����|'[з���!�vp�.�Y[�a��"��gf�����Z��<-�%>�{py4g�U��V3���+�#����(�4��D���Ø�ħd�JS�����p�8��cn ;6!�T`Q�ac�b��CZ�ڄ'C�`h�W�/��DŃ8=:K��Sc����g���u&QЂ"rj�֢�b_!
[�3��W'����$U˪�u|��S�/;6�saV�wy��1�ޞ�J�����b�ҳ�F��H�V����9���� f M�Q�{{���o4<AKP8���R�E��n}֣B|�g0��Va��F�����.Wg>=Y���7�b�ɼ�LY����\͂������,�|���9������ɠ���ӄ��z�~X���c�2�+L��[@���Γ��<�H��~O�ΑNj� �$>&�����F,�/�y4c���R���	��̕���k7i(	�+!EZ��jz��X�v���!1���4�����^��}[��/Lôˮ��!���]89�~T��(�mb�狋���o7�s�0�C�+�W� �x���L��k=Y7��Q���]?T8Ahn����(�����wx�:Ex�J����j�ֈ"eD���x=��w��ؐ^LE�m�9V���{U�
�7:m�������	��v�p��~�2*�\[�ƨd�M5��Q�ۑE����3	5�n�3��a�MG�T
�������{a��_�Q�[��%��a��mڷ[+�.�z{ ��+T�qǹ��ݽ���]r���N^fo/%����oc��H.���*7L�Y��/�F����^��$q�L�2u���S��k�[a�ؑ}?e��6�B7g{�x��8����em�����Tc�X%�^Y_�;z.�jKtLD8H�2�Ejb�
��ϰA��n�5^�ҒYXa��7(O��"�X�}�/���F�4�իf�UH#!���Y�,4>�C0�Q��l��=. �G�Z�D+4�ss ��ft�76�P޺ui'}��AJҏ����:����X.
#�����sP<�G*��w�~�B׳� i� _�;�6�\���`���t�%T���=����M<l�\��Q���~��>�-���@M��~(57��,u�?N����Z�A�d�3�]��C�h�n��|?��hQ�RP���	�M���Q�B!D$&[�¢����`9K��X�V�(�+���y��%��U?���������%�e�2E�jL�O���<?B���1|h]#`��]��P��!�5�Z4'�.�Ɲ(k�é3����m�w7��θ�:H��p{5���]ט%���U�[�����ex�b�e�R����lO	x��L�ːȰ>�驘/�
c�Q1�ep�5/�9	Z���njO�L�������"��2Qt��$�7^&	e�%U�= T�(m�K[�ȹ({&Ňf0���V��� �"��k��,!S�
��m}�وH���q	!�*�Qcn�0/߳�}hUo"�����:6k^U�},I�s�����O����J!��l3�EF�F%N�T�/M=0�����3��).�{����ˏ��/m(D��j�z�6M��B�V�My-����~�|��S�?�{(�Y���-������3��i+��n�,}�~:0�w�`E4U7��ˎF�����P�)1�6<�����Ԓz�]dR��_z�����>x��zJ���X�x�I��8R&���G>w:����΍�j�f�c;���Ks�_�1' кשR�r~	��\+�; ���&���H��+'�&��K�c�$X� Y�GP�LjE�U>T�YZ����͋�4�D'z�Kv@�U���/?*��L9h�������o�L�O2.�V9;��o]T^�/�
����n~x-\�� T�����,R�u��v�J!��$�kU�9��͎�����
�{����bvo��[J��-�S����~����hB���^4
K%4�Ø�~J�	���w��{Ƞ#N.������[�Hmiw�;�r�Fl�>Q1q#�>�{�Hat�����V&ξOQ4�"����9�;���5��os�$/�I�
�ǒ�x����`��*�m�4��`��������j�C��/��hY��ݛ���9��y�G�!	j0q���-"���6��Gl�|���<6��I�����	$;g�;�^�:iO�7��_���?�!#�7=X�$�_�F���,�㔒���p�/wDk��.�6��-:]�r����E�΅�X0�
0o�ķ~IN+��+L6S�T��%�|�J�^�moc������J��0�#���a�ȃ[#��x��A�M�J��1h����:my����=zbt��zq�B 6�Ly%��6�}�N��=�8��j��˺ݓ4>���m�,��.��8Cz��d���:4[�����Z�euX5,u@y���v�����I-iGuؒ��;��W�d��S#�r�9�##W�+Oc�T�Ce#9�W�ff޵=��9|NhH��=q�@"{��}�R0�b~�e/(N�j)DY�w�W���:Q�_e�?]k�7H&���
�b��@������̼+*o�ӵ@�)r������w���a�snd�Q��C���ݳ?�#�ܼ���WA;�#���WPS]�$:E���</ft�_������)_�00Ěu'�p.;��/ [�:S��<	�G�*��Qf[d�����3��j�41�~�`h��:i�y�J�~ٕ����6H���a�>��f�6�Kb"<(�<�O��d���Z���v	߄�~��t]Y9����E�w��$�������ZZ�%�{���tb����m׶��*�~�PX4��Þ��7 ��ik�6�s��MSn�c�*��,30�1)1�:�?R�J����.��G`"�����-��"�0����.�h��:Ep���g��V�#YlR�U}��&z���c�"��z{�̈́ٳ^���N�7mݩ!�ӄ�����f��k��Q�b��R��6}	'�eǢ��:C{;K�uu{��C��D:5��� ����A���Ժ7? ۞��ޢ���2l����>&��$�4b�v{��%��ɠ�����^�e�����l4�7�<�w�V����ft��]���FX9��T���%���p��=�فðJ��ğv��FqnCc���&2㡵�|E����z�=~G��2���A!]l��ۓ\�<#�/�yg�|�4�"fh`.rMPt��hy@259�}{�jb��̒��s�������҂������+@��rV|)��iR��?T<T�ѓ�u�D1hK�"�S!9&����~!)��!!�� d��� Y�q�0�d���_o�͟=$d�Q:Y�(IE�@�3Ô	���)�bg��v�{�d�م������ ��B����g���SB��*�]�1� ��L��w�G���f�=s�YLbJ&����v"�"H�I�n�3d�Ρy6 �X������������|�LC�i!��3��7�����5�L�	AAn���
t��u=K���s<V�~����/f���k���z�^��p[�2�;�� l3^���Ky���l��YH�ůV�<-��C�U���7$E��B.���i�(+
�μ���������I�Ș�'��w����ܫ���6�ԯ�Ƌ���"Z�Y�R�j�Yy�iRi�^�y5�[�=�R�>���er��^�瑓��J�.?j�*�l�}���*qn@Ba3���XJ�#_�<8���d���_ҍƔ����8ٲlĎ��Hzu���q�4���zbf�u�; Y5��;�Ay�N�	�B�F@!�!�5��v���K띚3L��|��-�r�}-�O�MS]�S�+{U�;�v�P�6��N��R-����%mE�� L��M��ԓgA�_%tӆn�`e9����ǚ��\����^��Z���L�Cq�x>3�qY�[1*���=��֒g��έ>B5������k�&0�E� I���+�P�ޔ���P���ѵ�U�����K _ى��y��(�'}��f�:t5QZ��a���beB�i��.�r�jpV�BK��¡B�ЦV9��+����]Fr#������|��;�/�qu7
y�Ŵ���Y܄���Ź���.�d���k�e��%�[G~{�ٮ�?0]�'�5p������-�%p]ī�%*���˽w��p��ip�RC����;���`<4u~�准���J�����#���)o��yN�B�L �I�"�����V}�VbO;%:�+M�[���jԎ	5�_&��M��y�!T��痢�&�qb�h4����uWSD�`���B��W��7����tML���liU��9yӹ�'�<��R�������]õK�/��ă��;�X��^۸���.�_sS��I�;�R]���B��^�h�-h{"�}�K����&v#� [Dm�O����c��oT�v� �c�u�vQb�K�(g=����S���Y0]�td�K�X	���/ИO+�X��|>��+x�YH�3@aeB�rhO!a����>FI�B�`�j���zh�@��ZUՁgT���d�i���{��F�٪�%�z=}Pã�b�F<X&�U�b�gu)�~8{1�����|����^���'@�f�-�pj،��Ԑ�v�<��<3��+KD��]B���������믌��{T7x�)_���T�?�#�L������U�d:I��!�z��t!�X���S����lU�I�3��c֣����i�zE
\M��� �Vk�&��ӡ�3d�m�ˊ8�,�mĶΔ�V�gwk��̋��V�����@�C|Z���h��"��V��6����Z(G3�T�,�C�:�K d{�n*ΰ%�|�� t#eV��ӯ�5���x��&C{VC�;�Q���eQ���@��a��6�n��w
��,��K��1�d��9����Sw��6~<�9|�ƋX_jT�� ��+&���ј��z��~��&���*]o�I�ߥ:��Q��<��z�$��gso�5�`��h�(V�g���g( �﮼�j���Q��qD�L�� 
�&�.���fd{��Dj�z�;�k�'7��/<y-в���I�%7���^O4���r�"����� .���\�e]�RC>�I�ӒG�讂.�[�i�<Jt���p[���s�����D3;�\�Dm?�2�di��6���*´��{���
����V����K��߆�8���8��C���Q�2�]��n=WQ���~�ȳ�#h���{cq2�{�����%���)0��/�۽2Qy��S��v�~^^���T��<�f��|ځ|������ ����%.aJv��0�)��-���
�E�!�y�)X��R �e����\��$e����"�]OOu�J���H����R\�7�/֗�b��r!vۣ%ƨA��۵l?��R��L[&
v�ga%.�Q6��aئl�����6��0��Y��XQwo1W
�a��;��* �Xo\��zn�KkN��L-����~&*�RB�-��)Ei3�ߙpYyB�F�Fi�������53������]�bhJu���~�_OB��-e�ۮz��H���$�$�kS!L���֩a�@��>�`�b'��`1��2�*p��� R���\�{u��JS�p�|���.�&����.�ǚjcx3E�4�Ɋ����a3�ЭUZ^A�qz�Y.�;	��vK���ϫ�D��S���W��\4��3z
���kWbr���WHj����:Cӛ�S���zM������E�Ӂ$�䊖�M��o������:��Hs������p�{� x�N�MB*�3,)CI?����F����IQK�8)<L4��.R�- bm����؛��𖼻�}0	�K�ۈFFƾJk���]���$����V��Et����V��Rg־�o�O?}"�U�
����E������� A�\r'(���y<�J�
�oGΔ3���G��U�Mv�Z �[�Ҽ���9�Ḏ���4ZY?��������ޥ�h6>��p1`m��Ce��X{c��-� G�ҙ��v�R���x�G��Y�)�D���ǟ����]l綬��[�r|c��������aG��&p�rq���#�֏��T.y���&�^�w����
O�|.x"�9�o'�2��e~y����,�XO@�ڵ
��X��-�!&S�� -�K"\�w;�-�P��l�}ep�3�B���Յ�]s�Ԗ�=U�O~��m+��D�X���a�3ʒ�^������e��ϥsB���j�����j9(j'�6�-��h�6�U�����=�cq�7�� �tX6ѿ��m(�i�ƃ�N�rR�|��rXR~���+�|ea=�f'���sK�uۧ�.m��挃"&�xN��/�������y�/����<D�Q|2�M$G�}��(t�W���S�d�t�mj�uo���n�K@ۧ��bk����m�Ooݽ�����ym`s|�"C6H�н��-V�qz��f���<�>��?0��=:I	�P��ejc��:�E�F�RT�C��L ��?L�)h��u���Q ��c���Z);��sG��F�hb&�F6��xpָ�o�4/kpa��ok�xl����	���.<�~U��4F�BB��%<9a �ʔ��_�Y=jQ�b��0>�����-崣�,�\�=�Y��x�L!, ��F��]��Jz�ۍ0�(=SC8��j���Zfʃ㪒r"2Va��>Q ��݋�]j��SF��X���0IU�fP����;�qXB=��\X�J�*m^z�L2W.�}eDDޖa1��wA���iMm�['7�Q�?��rxh�&�l�4�'*E�����1�:-�Z���c��k*�����/�X
.���Gk���B��݂ �� �ׄ�q��N���M����>�6[��D� �?��[z��}�PI/iy����j<�0m��̊O�ӊ�hV�h�84{M� lЛ뷳j�16�^��'	7����ΡWm.�nGyB��cɴ�ʎ����#��#�\.�6��F�:��}U>'�n-��@�P����=PS:��-�s
�f��L�H�cL�F]���w���7��@���4��簯�ȶ�6��)��H^�;s�����0��H�+z^C���}�T�qhd�qz�F�:T�#����WaN=&A���<C)���c�:�b�ҥ���sPb�`]Ң��M���2��/�yC������O
'�Н��HG���9���"�&ވ��͢l	��-����g�H��V�����<�@qRbMu���Nx��OӢz|5��c�chR����[�U�T��j���6�Mu?*j�{vʉ��,X�ǧ�~���6ukt��$�>J����2p4>�:����_3�5���Ư��f��ƾ��?x.U�4֣Y���@��ߋ���g �`<]��\����{�n�@���[F�ս�0V�
7hd�Up,��0	��G#��H�����M���t����:�I���UcyZr�O+_&�!@{B�Dքk��t�UXu[x����4����!(bb�4�u���&���e�?Ҟ�+�*ཾ�\Цn��Oe�Q#��6�i�X�T�NC�XZ��DZ�3>�$�e"YeZ�p������8WJ�d����mNnK�#w.�=/P��a5�F�?&4\��s��?=��ܾ��>�U�\��tP�?��ȷt�CĹ�ݔ!�.��gK��k ��{L�ٟ`�f�1��K�M�t���o�;��[��}���I�kE4����F�${��"�&������� ��ɯg{�qV���Ѣv;�w����ϭ��U��]�QH!�7��N��dӊI?����e��Kh���}��K�+�s����5��j(p���n��˵"h(��*i}��r����H���~Æ)�
������eGm�d���c�V��$�P��.łl����m[1���׆
X:�}F�L�$1��YwS �Q����})t�5K侂P��N鄁���E�!�<��<<le���p��Is�~V׷'2�\�5� u�
������m<L�W},5�V�j�+��s׸�Y���y��}���&ݛ�� bMr�Zz�w3'b���]���{Fa�js,ð�x1�u�>4OAtQ_Td�P��M�Φr�2v9�3����b���}�(۱}w- x-a�y����)��]����`qٚ�������,9�H54��Մ@�;evތ5<d>�ń��j[U�������z_��j��̣�߬4�~=�:����7���c�q�]S{���Q�9ځ���+C��w�Q�}� Q�"/���½=8K�(f�A�n]G5[�ԣ�9�a8̎��D졺F�ا�I��9}W(�;B��`��Kck:���	����I�}*8d�$�B�)�����s�ӧloIH��qs#�����)V=
�{]|��]�+^)���"@׵��Ѥ��1�����U����8�u��M�3��!�~?Mj�D�ѰC�Ϧ�N��T� oe*��E4z)���qA�:j�G�rL�;<7�fL⣈n�(w�Q�������j�u6���S-6���t�����ȟj�����X~B4@�8���LĦd�ͯ�I5Yfl]4ʏEJgk~}�j�OE'nT��H��	�Ĺ�	Cǵ$:<1E�g����5$2a%����$�5�y����F9&!�3��:{�>�]>5ғU��y�"s���x
�z���e�o��%�9��`���,� �����Ժ�H׊۠q
$����9\{ �!
�a�M.C�,nN���ʄN�6�Q*�#�He����P-fHrsB�B����䝼���9�_.a
^ 2	�&rk\¤I���ʀ�l3u��gX�g�XJ���*�������cG����t�q+��b6n���.���K�aUý�c����O�fC��k��>���a���'O
�`L��[B8~ln�n'�E��5Ff*����cs�p9<M�U(5-�-���+~B[�(%�����\X��v]�+�r�X��O;q����3-gp�&�!��V2�<"�2�ϸ�*�d1Y�-� q��Iv+$��U)�`��K���앢�N�t7斑�$���%%1;&؄��\]�Q_��8ߍ[�#���P��nӔ�+صQj����Y��w�ܸo>���Y��Ʃ�y�(�£%��b��9��*��v�`���Y��r��S^����Q�O*-�r�b�Y�cW������6#P�.e �����h�"+�~�H^��w����uU��-1�[��n>�&%�x�<�w�m��\��Z�����A�D��]�(���>FKʃ�J�H�4��UL>�@�E.�S_�u'Y�YQ�^g�qC�ho��q�|�|A�Px<��a�A�|��R�Jws�e(��4��Պgp�<���XZ��bD"Ŵ_;�z�k��ݑ�l��\!�T�x��N�_0���O���\��^�䩰��
��X�g���k9���Y��Gd�L+���W�2�ln6G�	�Jb�J�/Q��b�e�r���j��;E{�����Q~�LX�_��&>���L*/-k?���K����5�t!0�M��3��<���X�.��V��#3�0�,��X�j�.��^&Q����v��-�c��\q��oZף�lg���jBr/�s��ꈾ�0�� #3T+Ǚ�P��j�@��T���L��N�*��5!7�BuF�[�e��9��=�I���C72,18:uT�ɒ�[�Ah�b0�{�{N<5�D��=��=ȜO��@-B
�?=o�����<��/��Y_���=��v�_F�(�ib��z3Tv�����fdc�t�	 .�(�IrTv����N�{�D��Z/&����y��x��S��eeS��Ž!���v�P6^8d�o��ES���< <tK�T�Ό�o�����M8sp���������Bqm�$�$C4�p��hO�q�&�4����A c���?rC.ydrU)���8����Nz��Mϔ�-*���q}q�ү�9Ab*X�1�of��c�\�Y����M$+k�)0���R��~@��ܩ���HvD�o�;&�/��n�9��W��˖����=1Z�-�M��ؤ̫��י#�@���ҔoF�_!�Bf�z���RГ�5Oʒ�TvN����K���$�E]Y��Ii���Px|=$p�r���nUz��YM�*�Ғ��g=̺wk��L���!����"��PSU8�e ��L��5X�"6�4G�	y����-�,�&�K�K[ܸs���i���"���?~$y�Ud��i�*�\�+���v^3�C��Z���6��3Q� �C	v{'�%8(w����>6�����X���o)����r�ҵ�����\hD?��~t��OUA�T��*q$�`+ᐞO�ea�_1�ĸ2�~f��W6rO��M�C틦�"4���%l>9�?5/oŋ	2���"����68�R;�pN �d�ק��o3�s�m�i�׭D�*,���ae<ω��<�T�)��Ӡ����b�h�v�H�x���E9�J����K>,�k=�S�;��-h8xcmv����7}�I��|1�5T	�R��~�a���/�i� b0�m:ܚLnb75��U�0Cgg](��.� ;#4����I��y�a�~O���}��dvz2�����V˦2)���_?U�-�S�[8W���{��Z3��0F%���oЛ��CK���QP쑴^�!v�`��8��m6��19�s.�l�6��!(d*U����Gѩad5��:�������/:u%;�rq
�zIt#�&�V��cG���+ޠ>Fr��$2�G�06�&�ł�������٫&�#�w�=X\�MpjoYs��6�8���JO�s��S�X�2g'<f�ܳ�oL����e\|K.�7�vm�[af[ȥgl��6���,LjJ�R��5
���K�p)��>
Z~&9a��:)8��"���	X��*�Aa&�󅄠�νW��>��V~��;��L��.?�����s
���,ұ���!����M�z�И)X(��V��*��wS�
4�%��#���� [爠�.�h��AI�P���-���͸�I��5x`s|����V�me��cƢy�ͣ)�|�9<��C��<�w��]��ⴘ��yi��s�1U���^�	,��-�����G�1��>�����ߛ���)2_{�1.���X���1��M,�]�'�Bf��/�;�%����oF|���D��* �T�OG�Đ��V�X=\A�v1Nt�kB�s�H/&B±� �`sL�I�u��64Q'o��n&��?��2�-���%�8��q}���PU��lU�lV���N�����9^�����L���](���tCꠀ<7�����X�j�tߦ����F�U`���]'�l�@�$�r�(�6_�j���5�7�B��e���-QS%,o-�-�-#dzz�����$������/C�A��Y�3��׀��T��[�3��kx����h�A&j~�ƶ�+sH#
f(I(��G�ՃN��hH!��=`5L:�� �l;%�R��+�����X?L��}��Pv�����oBc�Va%.ەꩅbmj:bA�|{�o[�^�J��I�^�#�J�R�	N���:�6���d>�-߭yŊ��.B��<Ӗ��ĞQ@��_6��n���4Pk 庻����͛����հ�#{�b�H� m�޽�l�D�����K���
,�j�q��YZU��ٶBb{ً]m;n��*�w�q,^B���<�w)ϔ7�V�3|���na/����H-43}.6!�~γw�	�)L7�wa���:/v��1�� |I�p�˽!<ó:cV8;	qU8��$?�N�k|ْؔ�j��I�1׽��6
|�:MTK�M�8:޳T�?�H�{�y����ߢh�9>�k�z�ٕr�hQ�8Lv1�j��Mt<�[Bo����i�r�l|�Y�f��H�@��G-^�Ͷ
���f�_=�Z��Bfā�%xw���(�~7�][�,4h-���	/e�C*5��r��8A�֋�{�#ڭ|�#ϲ�k������Np0�3^}ϾQZ�L�*�6�5��)�#[�9�oM��:F,�4T3��؄���ۏ�Y���p��W��&�8���H�t3u9*�=�ҍ�\����_�������J̛T�2̏VΞ8FF0��'򒲊�P/E`=Cڟ821�Y��$��H����wl4�[�DQߟe��&�ae;�BCS�� ���3#E�P��uB5Ps�:穭�̨9:z��(T�8�������+0���Rͅ&VK�_� ��J���Z"yh8)�{.�2�,���\��M�ǯ�1�s����7�(3�vXv]�4|ܮ�o
��N;#M��y�I��(�C"��e.�¶>�U)�EJ�DW��Gn�h�(�f{��� �4JB�P��jr�eA���4���w���Ӱ�/��%;0��ER0 �`��v����pe���WPW���H�=�<A�����W��5�a��Ϙ��NU��{}�{�ZY�l�6�2�VM��.��~`_�C�cl�G�}�)��� ������`�l������V�n���A5�����<��/`�+�N(�b����"����/�Z��D�Q�V�X�&�&Y��쿈t:1�>�, y�	�}��{Ok�X���H��V'��F�,�͐Hp�B']>�-��Z<w��t��4�W*��xP��@�~�����6�)��j�4�e�V�KmZ������ U�c���kE�����{�ݘ����:Oܻ���O{�u#�G��!z�x{��aDRpSQ��rK`Z�� ��S�ޙu�~�xЁ��)��A������7����rB�Y/����A�B�X6�~��x&�-!�&�$<���_�[�
����|�U����|���#f$��%��RCQ��(BZ�p�*���d�gɫ���ڴK��5W�i�B �ۯ����үFs��~�p�<�o�����i����h//����<A���:������M�( ���J�"�ho���]'|M���I~$�Xو�Ӹ��ؐ��}{@��i׼�Υ&2a�b�[�q�a�0F1n�����s�ڨ20��� ��t���+ϙ�;o�g�W�+��g�/%�|��xՈ��������@1^��*Ɓ�DP��S	�����6􁡶+��m���Y�57��-"'CY�[�L4=a>:�B�$!xխ��=F�S񥪭
t�`�j*���A,��t5V�*]lDf�9.	Z��7���A��`���¤*5ml�,�D+�*���A��WDe%P�I��+��2���m�s�x	cz���9��DJ��� Ms[rN��G�"I����^l��G�� 3:~t	
��l��J:'�o�>��	��W�_�+m'������}��Q�f���|I���M��V�KЩ�:<��SӚE�F��m��u��Yh�v���{>���i@0"���3xމ��]��q-�y��-��eX	ر������|���K��`�ܾ��M�p�����[����	N�>�r?}��䨛�{�$%��Ж� b�m�%� �yH6PY��k��p5�I"�����g$տ��^�y9��\�I�$S"u��ǌ���B Y	�O�3�ի��8�Hώ��sTOcdrQ�Ut�W�ULȲ"����4�S�7 58I�������j�h��C?HP��J*[�F�QqEo���V�`���3k@$��"}9�����6��JP��.B�B�
��M� (�nF�͌�'��J���3V	�GO�bP96���Fv^
ҏ,Fw)jf�d��;��3�_�:y�X<��hg��G �=Y\mU�_�6}�7#L>^�'��f)�?��Y�Q��f��Z�o�����ɞ�t�j㖞�y���5����!=76B6*z�yԥIg�$��n�䆆�s{!�z�����$�+%aX�;`=p�zUѰ�C=�Y�
�#3���a�
-�8��<��=���r���`����eQ������edZ1 m�������8:#�j'�s�m�q�ꨰ�0���������C##Cr6o�߼@ٙ��)w���R��
~�hK:Mi�+���!�dC(T�|b��x��SB�����
�]���4���=͹#c�$�������F�h�iu("ȴ�A��!<�d�a��.�ǔ��*t���`�NɉM�s��M��3��;Sy�~��bL�5?ͯ���&�m�ͣ�@�R[h*�2P����Hɮ���p<Uq�r��TN�ޏQ��aT|�&~�;�qN�������r&��O�?���wTX�U^)G�L���grdt�[���7���j>�{�~�l[�"�T�-ӿ��@���*�f���9J�{�hg�|)�Lm��8v0������gc~��?�pBd�3�pM� �+!O��Ҝ��y[�I��v$5]���M��)����,X�x�ӟ"V��bƓ�DT��8��h�r�,�����J�x��vY�j`�|2`{W�Y�
�m
���҆Wq	���K'[�V�ҥ�Ũ��N�N�t0a���]����ʚj�1n�ss{I1q;:�������G��i5>Y�)`�2�gbOP�x(Pɶ�1Xo�.�s�S��=I0м��tm.��^��[�6y���T`�c�9Vh�@k����0I��pa�����V�9e�� c*;�A���� xl<ԩ�\�5�:����EN��E�Vja�K�U���w���V`��v+Ы$O	����ڿ��ӑ)
�c��X�gh�f��ŕ"'���S[���#�R�C���g`�d����#mM�>5O��Xb��d]�;�}�2���������k$�+�Rܔk��'h�v����9���$ffH�-��l�¥��
���U+M_c����L#g̥:�{F�j�d���k���g��1���ܨj����]�NZxR�0r /T������ƒ��C�N�nn2]n2Z��{�p�D�k��,s�e>ݰ���'fH0�B4	��k� `�Ӹ!F�Su�ȩ4��Q�r��U�k���%��dJ�֕��17؄���<;\Q��np�ٿ\H0b��?ӌ��K�|��AL�>�#�PW�E�؝P��;�Ԗ~/+Hz���v|�ZU�['�J��+��/�L��Q`P����vǖ�i���j:S5��n�¹�9-a�m�>���"R��ZHzX�(E���5	HK�J�N��M�.�L!g��S���QJ�Եj��\Y���vJ�]��_:�.˥��I��?DG�.��ɓ7��Q�����;l �y����n�ڡ��&�߶r����X��Z��rf�E�->��OF}��N�--���^�N41 ��#c����E����%x^ßL��h��Q8-%6u�6g��g��zI>ydy��M?k17|ҽz��u��ae��H��Sm�;(7݊zLqA�1�7F�@!��9�g�߫��ټܪӋ��4+ ��ݓ�� ��\B1�?��Zn�qCX�;��������nq\������6� g��E���S9l�3��K�Noq��S4Q��!�0Tզ�����)/]�4/�T�!���Jy�(44J�[�{C&����2��:ۙ�P1�B7�su����c�?0
̋�E���-�uM�8�p��*$�cԨ爕YG��LB�;5(�sJ4�/ �o��#2��b��.t�wQ�G�bX�8a���b*}c�&I��*洙������B
��9��F���l~y�>�2��A�/��[� �w��*��zSi�d�x��_��)�:�B{&�F�vg�0�?�~C�-�J�Y����Z%Xʬ��]��
�Z�7��Ҭs�dU����HT;I���#�^���	(O����!�A�T$�Kh �=%H��g"�k���1;�y��_��Rq�V�����&��tM/�/��Q�\xf���*���:2��q٪]����e|I0�E@�s�W=g���esU1x0DSS��7��H��:���l�BO��i#<�D�y'�ϻѻڧ�s^���K��4�R���"ǃoũ5{?@FZ��eAy�9YwE�\�U �CJF{�u�����M�������_KE�!�#
`k���Լ�g��^ݬ%*�¥�ߔ\�ꔓݐ��-
G� ���E�
o%��&UY��`}�/�m��s�r���F<��(�"8���ᐑ*�l�^%��N��=��%DsuD��4�]ATZ[�y��C�7����W�]U݂��0(^vO��/~wѳ�G�p�*���#u�?c�F���7�rD"�GG��ƥ�x�k�I�r�)�n+*���Cك�7n�Fhi7�̋KFc���ǐS��4	�G�'�r�O��7��˦B�kX���Ɵ��s�@�`Z�Kx��z�����v�kq��n1U@�<�׌v|�/O;^A���b�����:2���@�^�:��#��Q0-���if������m��������S�jY�F�����1,l.�:.ؓ��2��"�"�[ڰ1c(��>��(?��<�k>w�!�mqu��1U����KF�g��̊��t��-��(6B��7}Iq��{ʐko�u�X:��Ŗ��k�M���{ǠHWE%u���b^�ݣ9�Ϗ�T��&x�)K:�}�G��2�:��L�-��O�t��3��1rm,�a5�����2,J���s��+Nx���J�x�š^wj� �+]A-��!KHt"�,Y@@jS^��yO-qV��(�����ᶛ42��=�'c�����(���p��_6eܣ��V���4l#�:Y��cq����ځGT��4mv�%����y=�ۃ�Z��.�.��|�>�v���@m�ʸ��z���:�|	����B��������X�bzofUWNrv��W��Z�y2��׷��~�Ύ�u!�cj���<�C�;�w�hqleïo0#�Ζp m���tO�nU+p�M_z�whXC�;��.��1�ɯ��T��&�9E���n	jO�VФ��K�=�cOaJ��&��sLfNϽ�Xݽ��i��-�/.�P�"b�����#7ؒ,M������M!�*Z���m�h@��`R�iW�%�"Mq�6=�S���y��?�[�ǋw8O�P_MdRJ���R䇉��&IpN���+.�*ABdQx২��r��8�F����&>�Ƒ5�jP�~��T)�˼�dT����l��uU]BN~�lP�j����bfc�!*\_�n��(���Z���N���p�>��Ԧ�4��Q�@.ɄܕeG�85jc7�>��P�t�v��K/�|N%�߭���J���{J4�<���舋�^"SM���іߵ$�)5*����1�,J�q�"4��rnT�<^�	R!��b��{�%�@C��b�5�n��oJ^�-��&O��� ��-h���
�W���	�����jM�f*��8G���Ѡˆ�t��������R��g���8:JU� ��5�O�Q�z�@�{�����/��Q3\�G�����ȣ�:��]�r�[�"��]�05���X���3�cȷ%����=��Zl|�S}�e���n�q�V��B�K��X���42������S�7(�� e�k��T�ܦ?�K�b}7�;����]B�tvv�7��q�bcKb�e�l!�ҏ�l %��'� `������G��z����[��e>����(������.N�@%h�
6p2$*O��?�
V��+�KUjǁ������-��he�ĳ��F�\�����ld����T�G�w_����(3ġ1��!��T��I���}̡G�N��d���J
�+\Ωm���qI�D҆K�ǣ�{v��@�lU1�U"R�,��ZNgS��g���zK���������i��;�!82�u�pkЗ׭��NmH�p�J�5wƼ�";T$����6�2���~�/ٲ�<x��Y�Sy�Z�;2.X.?G��6P�.k��8]r�y蠰	�ڨ�,��^��p�:��\σ���Y��<�3e��L	�{8�l@��*�U]�W�H���T�R��κF�=��_k��e\m��sb�A�g"�<eqʯ)U��V&������_8���x
�iwiN_�]��x=`C�]\��?�H֍��d�Y��1ݝ�8��E���- F����L���D8�@T��by"�?Boj��1w��c,61��[H{\'���3��B�8�]d�}���D��;ت6���2��������,���w ��������W*���}QH0�׈�G����!�;>�f>���{����f��b/J���s6�k�V��{
j��r6��Ƈ7V�}i0�ӻހ�P,�#E�UM�X&A'0�pwJL>�D��)�h�2G<m��,��>���9;K�}_*�?>`�3���s�"�y�2�N���T	��x#�4��jI�܃2��3�1%�N��/t�O���T8^�PK�m~C�b���=e�(�"8�A;v�G||���|s�(�|�J��@�	��ʪ�U�nK�=���ݵ6��?D��G~�)܄�J�+R�	 �ԫ�����I�L0q��ݙ��e`�H	�m3Ѡ?T�����3O�Z\z�_�%o�S�>��^�	URO|2�|x>{!9W�f�.B�D�QW�s�A��ӕDh.f�m��L�R� c:Y�j\~c���(�fZ��4�%��N���������y�4�KcJ_q�p�L�9��:�y,����u&w?�[
@3B���n\-dD���R`[h*+k����#�ʆ{�I���a�@�/��y����D��DsƘ�d����r|��A:���c)w�,��}N�(e�i\��&������f��ύ�B?�ZxU��-�*,������%YF!ü����F���N�z�~v�sdU��~��c�jred�P��),�]�ϐ�83ٯ�|a3��9W���E�@�|��Ě�<�>Z��Ӽ<F8}����d$�X��[��9�n�9��\�g}#�ƮN����DV��6s�A���7��|�+4�/��6�L��U ��P��̓��O�L	�K&]��Gl�i�,�a4��tV5R<�Vq�3�(Z�O���L�V��G�'8Kp���nk0S���/9oZ]&R�������bf��L}>�d;�<�'$h�.(������������/�H�ｶ�
Z]Ĥ*���-����V$�\���p�Ri��8�P��'r�޲����?Ѵk�c�!~~���lxwx���WBd���m�����؝3�a�,������.��ܜ�.d��[y��M��g�>�\5�ð�(�gz)GDq��/o=�3J�/MU�����/%�?�6�)�c�\�J!���g�]���K_f�
��z�y�������x���������x�m����ܮm&?��n�[�Ͽ������]����Q-����Z�����$/�WN?�حz�"��՛�is�򵕧n�M��� t��'��6���(P�D���U_n<QH�Vдu���k�t6yw�62ᣴ����)C�'L>����&?l.�F;q*c�t�6e~P���]�
>��H�-:Z����y1���٩#Z��/�H�a�;��Rq���K<^yz�[i|T� !$���7�7��4ٮ��mT����.�g��L�A�=�Q�#�<<�]�w]8�����ʉk`����40����t>?R�<�d
�Y~�G���spt�|��{m�33��.'��5{n��D����t��}lH>�oU�� ���B}M3�nV�e_�ߘ�q�G�^������U��U,���Tڊ} �k� o���
GK4�\
��<�}�����U�=vʝ�2t�Uɭ�؟'�,V���.���+�5�OV
o; ���)i9� K�G&"u�� ��	2Vj�kJ��-��e�F�ӌ�`t��ySy	>���>r* 7�λC���[� ���D�E,B����0�L���|@��ӑh�z�m�{�Nbà��ޟB|�FH��g��H����U�_���=إa�;(����[����Y�KR{c��c����84����h�p'���b)j� �<�4���*�*7�,`�Zkn��݇
/W-E�RmTE�	i�k^p,�Ҿʉ�|���y��hg)v��˂�ekU�ݖ��v����U�,��[L/2�*ڼ�G��2�!G@]����s�ٻΖ���[�<e�Ÿ9�N�;[��B�e���b��݂�������BZ�8h~�xƑԠK�c���77�W���G�آ�
�ӧ�ǡG�m���g�݀��.��+�.�.��+E��]<0�&�T�z�\C; <k�9�I1!��]H��]�r6���^_�sghX�E��/G'5wM���@W˭�4!>�����x�;��x�>}#o�#)eR�2���'u�T��Y2��L����i�6�-� L�0L��&���Λ]���
�s@d��:w�{�
r�'�����"�9U9�IVuy�b�Z��
�q�|sf:{3��`&f'y�����:���̃���ʈ1�!��`���	*��҃6ʋ$�����o�m)�Q��5�4a
��۶*�4{�Y���o�a��8$8k�A��xu��X�v�HW+��1��u\ѫ��`��xZ|z�x �ա���2�{@��%�*x�k��<�.����r*ߙ��ǋ.��#�׬j��%]c�\~�<+��U:�����o��K�M(/0��;בY�GԲ�[/�]�K�tl�غ�?�!��G�Ճ���y��}�=��ѣidbӚ{�R'�Aet"�S�PwYn%�h�F�=��qz�K	mN�XM?
3�C��rq	oF#���(oC�:w��_�z_��k��J�@����~���4<��׏wg�,��/����&N�]����*�����ޒ����:)�����7�_��n���bx�m�����J�(��%��)���o�C��)7�i_�5�bS|����&�$Ý�&��G�3�e����H(�/z�T�Ѿ�M9���qB2Δ^vI۬��%�=����5,���+�Ȧs�F�a(��8W~Z�,3O|C��$�=f�A�-�Me�q�,��%��2����H�o��X89��b���Y%�Wæ���EE��c�aM�N�v�ޝPh0*뼥��&�vj���a%���<'���/��� �/�T��a����6��"���<��$���vC)��v<]��_X����kL�/5�nS9��]Y>�x���,�����0�P�׽��!�V����+����*��
Xy5�k)�I�B��Ƽ��o���B��)��K�xU��Q}��L�X��ܰ
���t������L�g=�C�W�vWW����}yj�_f���(���hgٹ������ށ]�`'�³u]ؔA;=��vV�IE�wc����m+0	������mB~��$s�%JMZ���Ge;��?|�H�Fr��`����wҁ��`��L�)�Qî����{^$�s�0c)ʡ2K�.#6�N��ؙe����'1�^H�C�C��LL�ց��^9;��y80�@w���\ї4^io���z
�&��
��#�ƙ�d�?~PQ���EN�鸤4��D:�h:er���a� �ܡ�ը��v�P��G����~�t���\l�����!�Q!y�{��c�r�o|"��� 4A+�w���+j1�"�9�O`��a���ƽ��Z����htz>Ć6�5��}�R����#�7u@~��.\���3�پZD�����5�:���a�hD3�,��w�l�M�gd\d��C��q�}�Y��%��:��w�sNC�o��+�Rؿ\޿���.i�L�U�u"#�D�n�(�;N���T!4��k��VuzR����� ����d�	��S�mb��9/����W4)-�@�-�P�;y`��?r�j�w�Ì �,�9^�gwaD3�K'a�z2�jң��Q�3'��(�֊���
�kn�ǉ������|ް��s��o��XC�rz.��Z��]����QD��aX2��Ut���숮 2e�"����(|SB9�*�ywDHv�ce#]��y�QS���+����ޥQq`~���=�:�*F9��i���r�X�����k5
�G�@x���ԛҀ.�s���{�3�"��U�����i��s��VW>��V�`���}0�(��i��m|#c����Q�5��T(��&�H���#گ+��W�������m4�����/V>6��R�Y�3/L��}/�(��YdE��B�U�ِ30�P�����3(I2��#����j�l����]}D���;���u<�<�����=�N�Z� ��>�^�(�lt�[+�7K�̺���
~Ia/�3b� �0�4����y�}�bʛKޜ��`���n���=
9}kS�5����T`cU˦u����DA�;�]�4���a5
�W�:~�V�(�)$EO��/�cq
z��;Q���G;�c��B �	;3�NҖ�)kЮ�p��Էعfۛ�����l?��{K����I��X���fh&hR���u�{-�Zʑ�+��1a!W�KPI!�6m#�'_׹��`���
<E)<�;�hB(?8�&(ܘ@�!QBg�z��<�����]=�7������{ b�����"��~:���v&3O�2i�W��z6�8���P,q=Ma9=�2?n@!F��Ҫ�IE;�Y�X���Y�l��	���q-J���������m�U/�@"ΎO
��Y��r�n/	c��"|+ #�CJ���G9N����T6� *7���<SH�hJ{��4��f/�oAY�.�q�"������O�G�H��>�t�g˴��B��:�2B@VMX��zn�ګ�o��Ҁ}����$����I�,���6E��攉})r�y�t�s{/��D�7�m��U/��\��<BpI�P�����?����u?zQv�4+:�b�o���bݍ�@��	:(��V��`��S�Έ�2AOeg��by-�vK9�^WH��Q&��\J^b�PD?P��"�b�+�c܀]GR�`��P^
rW�G�u��
[��B�;E�ex������5<?Ӳ�?�"�euJ�k
i�H߸�_���j����B���� �}DLw\��C�SLe�٘^h1xݕP9��S�:�Ƈ6W��9�y�+�Il�K
��$1/Ez�r��#�g�8�(����k3�7�n��ٝ��t�d�K�8�w�H~���_}���3d��l���I`ca��t�������UK�q�OV�]�T���`/���'���^Ol(6z Brӹ�ڱ8�Lĕ���$n�b�W]R��ԂZ恄��ӽs�B����9gYk�?�!R	PZN����b�
�,|k��m����}�I���m�0�_��Ao/�J�bz�ICmF��a���I�p�Q�u�]P�I_zTl�����v��sn��g�k̶��}���
�g"�n�mI��濳��~�S��� ���YDQV���L�V�T�a��幓�jH&ݞ��K����)y�����8�X��=�S����Q_-2��\�gg�W�u��}�S��&;!]^rX�-�Qʡ�'x�	]-��tB'�bt�a�V�v�+�7b̒Ȑkj]���щ+�lB����`͎�[��dW�u�}r�m�i��La��A��-�Sܚ����!魹�bo�{�B>pQ�!T����0!��zآ�aH.�	�����"*;�vہ����?6���p��N����UU ܈�߷�ǴQ�������r�����=�~��!��R#��Ӏ+�X�;��e*�$�/�M���B�\�	���<���^�V������Ym�~Ufy���ٶ�
�[�D!]:E�鑭����E��Yz��љR=)�]���7�WJ�5�Ԯ�H��E�e��g�BbP`��`=�(���X>��y�Łd`�C�-e�.@�>i[�
��{��I+�����3���7n�!�V|6@nmS�⛯L��p,;�L�NK�v�����83�C�p_�FY.���^)�K��A�A�/~�c�\�O�g�;��r>�㶕X��go��ҽ� YY�O�ξqh�-��$;�iy�Y�/,PD�U�C���q�]V�㰠�ؼE�Q�T�W�z�1�}�V�[y�2 濻K]�s��=��9e,=��Z���b���߿��h)�����(��"�s:�h�m7��9��{�?�K���L �xpa?{���oe�S�l��B���b|��H�0+]ت��Y8,��q�+y)�ER�>(�'.��ksYY5���Et|���}�7U<���\w6��� �䁃/Q�V흢��
�7b�b1�&N�����O;�/��LuNͤ;j�����8�ɐ�j�8%T��ĄO�L�i����
��IbV�����h�C�ց�.C*(�:��!�Eg����F�RQC�M�K"�v�a���<�TC�:d���%F�a.%�йT��.��#�!1ya�@E�k6��ـ���J����i������mgj''��[ǝi8
1y�F�=�k^�a\���#Gzo��H6}ڭ6 �)����A��F֚���_�p�J�]|�����B�$�4�۾t�H�Q=�s@�.7�= ��PE�;�4^iԉA���&ҥ��������W���]��~��׏+����	�=2
�S��߬�����Q�xs4+�:��+f�7v�#*AW��1��ԁ����<N3AUv�~�i:r�
b��=�n�D�,c��)�k������=�C�`=�Mo~��s�	�7��ަ�!�U�f^��D�����ו�$}?�Y���Hv�$�i��ݤbxB�ӗ���,�`�����0��j�J_�>
��8D}2�cN��;�u$c��\�R@8�4)8^�1�2�+�r�֏I��nV��Aܗ(,2���`0?�.�'ژ�V�C����^�߰A��qW�A>�-�� �?��S�?�
l��O���z��ǘ�;�����;���x�zm����p`ee�s����^�pf�X���33a3�V��a�8S���ةJֱ<� ���aO��و�e]�'���˥�qs��ʌ����/A^�N�H{�!��CdQ]�}J����	``�4�:NS�5�-jW�	���,�N��V����A������w'uV֍/�5xUf9�p\�ڇ�s�t;�&��9;��O �
��Bx����w��v��u .d_<���oH�unݿ��ۅ�3�c��Ǝ ����vL�_��褋�C=,����v�&�T�S��p�!h8��5���&�0!��h�!�o)+���$�7�eTiPB���V���C[��!�zj��8�@8HO�Jz�C&�5����6�8���:YSB�V��N<�O���k56��qrn_��F��˵��y9x�9��yv���jYu`E���͓T��RM��gL1�[�G�ڿ�xK��qX��_�Hhv�P��
��"��+�~��X֌�����u����
ԕ:c��`�it�<�)�W:L�g!"��{�?
Z`@�F[���H5e��"~�Œ�X���]����-8�s)�bʔjJ��3�x��e���c���3�ǈ��������qcz�U�w��%�<_
+>�p$�0���:����x�����z�y^�!_�Ir"��"�̅�pȁ�fᷕ�`Q!ANdCi�ҁ��w��ZY9"d6�W������?��D�~���f��G^�o� �L@��}��ќ������O��sO���:���e��!�7X�|R�$,@[g��0bs$UOU���52sB_�#�ӿʅ~��*0��'�H)�\�p#@���ݥ���~��M����@e�@��6�m7�}#w OC3��"�h� �o�J�����Mq�2����b^��*�<*���w4ף���o��j�:7�{��;2�c���������)6A��!o�h�����D��
E�]r\�|�Z|	M�6�~d���X���iI���8kA�סS�������K'�1����Hc���Zp8�ұ��s��x��Ӱ�D�FiO�@�A<�.e6L�iGX|i�ұ�Wѧ�q�B��������b�}�m���l�L�A���Sz#q�;z����p�5'-eцMO6&�����j#���t�2��e����1����H0�.�CKU'�6��c�{�o��A�T�K��"�ڐo�P��a������xU��T�Sa��E?��g�q���I�:�!o�];+&�D^��H �?�G�\w^�=*q����k޴���
�[�u�z��\�uͳ������f'g~��,*�9������2E!C�!|	�3��g��-r���"�Ö
H�o�#L53�
[�rNK�r����Ѭ�)�n��=J	|5�;���;�ݜk���v�%b{z����uUfՑ��u��9�L�rM'	�M>�Ȉ��h�1���S����/�b`�[��|"�I&@��-�~n��aV��9�=����%��C���dL��U�#�M������+��[�>g�!Vx��|��|2}/�B)ͳ���Vu}����@_�VHe����ͅ7��_J�#u3��gq�R���f�?��q����~�4�=d�Wr���搌���g����:�KM�����0�Ě'��og����8[����MIZ�þ��e�5,/bɤӥ?����$����Oy��b?*�;&"S��M@ܤ�A:etB=ނ��x�TݡlcC-W�����{H�B��#���+�E`�f���Ԣ;ău����c�g�7*Ee�.o�y��fzG��mI�U�~č-7�����+���bo(KJ\5B{*J��P$8��gH��~�l�wB��a��y�Q��\r�Ey�C.Qª�z*���Z¨����ul(�I�F�Y8Vx�dwJ_��Ҧ8��At��\:�i�,<m"���W���Ҡ�G6K�hbPfǕ�E�Y��+�r��Г� ɗG��I��i�o%�^s
�r�pz_s�9-����� ���Ѷj!���8�e������q����Q�`��߮I�C��x4���C��?�G0��O[�F2c"��1l�<�<>�Ӫ1T;���i~GÀ"}����H�����%Z��yW�gx���Q����eq��qzK2z�S��Ցʦ.�Ny��'��{����,.Q�,�q�vE��E%�$idحB���1�( �T��i#�Qq�1�� ���.�ޘ�p,�����f�_�W�w�v7H�Z�,��Ʀ��L��b;���X|���T�sp�q�����G���?t��Й��;md(WY��-���*�G��,a?��}l�h"}��ۘ��f}'��w�sC �tmh@����#2�-�����C��Y�:���N#T`���%��-0+�G��2��V�l�_�*�hM�Z��©H�F��� �1ح$_�:o��4�g-��+��Ա��v���̖}vJ���7�l:�%<L2�3Q�f,K���أ� �+Q¢�b��X-1���s:5`(����cHk�t� ��_���q�iL"�m�xG�AP�R1��E��X�$��;)Վ�b� �x+m,_)#�t���h�@8��m��������ۤ�����T�%4[��H�(��9ߩJ� C����!��6���@�%_Z��0i�����w�̋�����Jx��IW�N|"�~�DvA�ԇ[D�.vCd���<� ���jFh�X�}1�k��,�-5��4��k��9��R�9�X[y�?��CPx(����b���;V�����n5��j>�W�\��9k���'hSz_�-��՟�q�)�͡�[l%�$��ܒY��Ϭ�aM��D�x47��k��^-j>��w�L1�:�YTa��F0`7$$<�b��I�?�|���ɤ��㐂����Y�cږ�$�G��Z/��������v�d˥0:�����D*�����>w6����/J��h�s�ih�?�m&=t9�H^nd�Z�1@=tr��i��ೡk�V��w�>�>?�A���n�R�D�"����A t��lX~hk���, Rz#�>#�Xz���pej:�镩�W�{�ɘ�rF.4�c4�e/c��hE���u5���h#��4�[!����A��P�lKX�W���g�L)*4̘�w͂��S�L�<�n� x���ӣ��O�]����D�<c�#��}4�]���.
��VHWor��e"� ��R�O��p#�NX,ԛ��j�\�i�"1�nC�ς�E��ܥ��e��#k�� �$h��hQ�ޑ�Sk
 ��s�i���.P�>���Q�#O�i^o���{%e�	�t�Z܃�j,�q}����U#+��԰��F;���zOʐL"�79}2ND���!��J��E)�TR�s T��J�@o��G��gA���i�2V����[�A���,>I���:�LbPu/
���e>�#�>�#��]w����ɳu؍~*{������̑�����$��ʹ?������'��F�:m,/,��(�<�Y�iV3�,=�+�C�m��)l
Ȳ����[�dn*��]�x��0_�����u/50�|w�̶�<R���չ�v�y�����*|T)���Y��u�o������<M��&�Sg��|8����:K�<�r�=J�Xk~&��ʗ����Ҍ31"e����l�!�� �?����|�/rp�#w�#pJYR�_ WH�G�j��q�gz������.kwGSs9��R��
�0'�Y�Nkq���(Cw��!�:-Q�^�Č�]ڐ.>Hf��Aڞ��-O��Z�&��[�Ab,� ���z�����x��4�B�c�����f�C��0%E0�p+A���4K��3�����N��&���gU�� ��Ho�^W��kx���2I��r�i'V�Ty8{E�n?:�c�j���I{���+��%�ZWȻ\�<�MJUW�Nd,9��B���l#�����&�:�� gC�d��#�����(�H���a�Ej#v�a��j�}$��B����{����>���ա����ý&X���΢C8��S;���_��9LX�o�s�y�I`+Ը�U�Zsv9{mr�COx���"��Fׄ^`"�
��Jom���k�κy�����	�� y�
��t�>!��^M�æ��n��LJ+kP 0o��H~B���i�h�W�M)�Bҭ���3Ʊ_�H�Д�[�{��Y�[�x��X˱ݏ�RK�=��y_�' O�:Q�0�IzV�y|�- �VYꉢ��A������_$!����_*q\<>@}/J8$��88�N���:���ƦD�CK�r����d�G\CJ&�Gtl���D�5T{�S7;N���V��&C��ckO�����'�&ޱV�CK��ݺV�"�����q����'�x'���)>��BԺ�'�u'�y'��{�TJ�W�����f(+8�����űNφ�������L�[.w��ֵ��
�~���@��.����L83���⃬����X�d�Z��a���f�xHZny� �פ6��1�b@o�ځ**^S͜��X"A�q����/��^:x_1ѯ���[�@g?*�	������Z��
נU@�w�1����V��H�"���,q�2�G���X�&�<-�1s\�����P3?<�.����ܼ���RО����͑T���tg����a�ݻ~������5fq�S�������l����r�����WTai�x��:i��ڔ@��I�#�Db7�h:m\\M����F��eAcfnK?��O�X���Rz���E��T�JZ�z�i@�k��n��qOP%��=ɷ�E�һ�U�5hz���g2f%�L�l���0+�����	'�"�&!�伌l�#�-�H
��Xx�Wz2���l���WZbe����-�j���`[#\�C8n2�<72�%��"�䗖9��1��iz|����n%����̓{�E�.���"!��ܺ� *�
��a�a����P(�f�o�=q�[���n�(��I�n��s��LJ�pc�E��B��-�ig���B=���~*fr��	�U38�=����T��w���q���NZ��_1�����N� C[�P��r�a>��[�H!�Tt��3lk�yɄ}�r��o)�p��6���bx�K��j8�''�с�͌��\���zE���o���E\Ϡ=��=�Y�bƗ���FE�3��j���ʪ���dzJ�9�O�=7��,j�:��^vSlE���"���M�f!����
� hC�̓���ѡ!;Q5<�B���G���S ��b�4����H�r���3�	�	E�9�.��k\����|��A�uj��'�*�&������kDq��a���ر(������L���G����� ����7�- ך_� �v��a	�S,޽R���z?4"��5>$���c�d�L�CO���$:�+|�U��L���r3r�r�r�c϶2�S;RZ�i.��1(�*�m�j�F���
ܐ���.����_͵���8��w�H�\u?6�X���=+�"���Y�'ﭛ�W�� g����0J72��I@y��JƂH�H��+�d��~��{��a*PY�k!9!{?ZR%��E�귿�������P�j���~� '6���mٓ�hSyts����(���4f��(\�p�z| d1F��#AU����e���U�vw�&�ە�+.��2ފ��|G]�N�r(�)QG�
�=�)G�t5�q�'�N��u�(EU�H)l��!(���Pt	[�YN�P��r�3O��g�C�p���^��L�o�0ijW(D`]i{�čۃ0�LF��� ��14�t�Y+���y!�]������`�X�Ë. xWF]A8��?=����'y�8�5��&�<=���u!��K��A]p�0f��
�#?O
��eد��"ދ�1$P)i�m-�������A������_�x��q��7�O�oM�-�p�C���44�yy���t�)s�`�
�o|�=7�/�h1�Sr2�EP��=��Ԣ��5�$���seO?�� ���g`j=�!���r�����V'�"�/����je&و#k��peal�Y �u�vk+��6}h+˞/��:6��Z�΂�lh�I(������!��4����@�K�:쨒v��D*�+�R��R�؜s:�&dw�Z;Y�:�� e���͙-��	�)Cr{'hǏ6�X�u�[@É���.�J�/˃�"�Z"�1y���y�"U��N����VW1h�Y�tO�T�C�Ɔ0K�C��O��O��;ۇJ���kK;��>O��E��6 ��]Q: D��*��+�K�xՎ&�S����#NVJ�.2���-����s`�=�$��`p?&#�&���� ����1�-��)��&�s�@iM1Aq�;�8=�~QQ�n#ċ��f����_�i��q�]>�(9�C�Y����vhp��YG�%���ʀW���?�z��?*�5�Xݘ7'���1�J�ܣ�i��4JH��Foo]X�.���^*�%�w�@�oj
	�A�D2)���K�[��N[������r��M妽����֝
�Gj���$N�:���9|\sz	!��U��B~8*�<g���62/����V��-l濇�k�^����Հ7�e�L�X��n����p�8B���)�r��5��\��ڤ��o��qK�U����4G-oqakY5`��fY��͹��@�0'}�Z���ExW�i{��g�Vuӈϡ��+z/,�?�0=��	Zt��!!��Te%ۄF;,J=WqY,M���\U�c5�\���� �0�wHxVLA7P.��7��7�eb�����_���q8�\��&g���,ڷZ�U�~�I��sœbԏ��N3��eX�3��K���_1t���>fQUZ�OqK����#Ũ5W��Y�٬�M g��yE��V74�01~��H�Fy0�o#�+dR��XI)�a�6}��%�5DPR��St��`8���4�Pc ��+`l�K��(��K���9�-u�5�O�n��=>̍}x D/em�cH\p�'� ,��T!Sܷz6�͉�ʪ�9X�1XT��D���	Y��P�ڴWğ������⿯�ƶ��C�ƹzm5Z�aH����W=!�]��&�#�VD����k*�#�VvG�F�
�v��ͩDnY9��p{KA,��1_����?�9�ӏ���Z)������K=u����|A'�*�~*������.�聢�c�Xk�A*��}����SY�,�+��cw_pm���W������R~���/b�`F�4Gn����S��,	�Nm_	\"[Q�g��������ւ��Ԝw�\���`��6f�?���UA��Eo��H��⫪=4�����d�k!�Q?�9 ��F綻�g#�,D�x,���B�=;����Z2�w^w�t�� (�
��z��>3�j^� Zc�83(�'�C�ج҃Y�nߦ�$1��_~��rC�kK�>�VL�7=�*�.O��]Sg���(�ebD�-��D���cx�i+{��-������WJ%��N��a�?`Ǩ K*��,B��������|h���TH�oF_����_<B[n��a/>��V�rPa��/�~��}��>A���N��e'%NH��\K�:2��S^���$l���#x9�<��-k�]�N-df�О0p��`���V��w<Nt����ƑD���@lȝ�U�b�uo�0B6e_l��з`B�0p��ȧẄ��݋=Ԏ5����b,�����.� C��L6�%�U����������M�9��m�yk��z�t�Z<1��<Z$s2y�Y,�u�e��������r�պ�i��Ԥ���ENoX�z)o�� �5�!+��b�^kS'���64ϱ?��-�#H>�U��c��h����I��#��>�[H�����
-�#��S蜆i$�a����A�`:7����ԙ!��jV&�_iu}q�v����Y�RáO5ښ<�����rb\����߻xC@��eiM��S�>ٶ8+�V88f�_�����d���og��W��sZj.ṰH�%;M��!)9�F��O�h[���²J�+%)�it��5�W{����"Y%	��TLԼ�ח
���9���#�z��;�&n�~h�X��@��@4�c^�H�����~���x�L�ל��3nӳ�V�N��5����xv���Q�2zE�Qا>�K9��9�{��/m���{Vo�Z�ѣ� �`���ML���#A�	�A<h[?}��79
����/��>"F���,'��
8y�a�&c#�>GW8AL)N���k��И��e"���O���8A��9��~
����P�11��2�%SE�*�6 ��!�ǥ�7�Y-l/'C(}G|�� �60�~s��,�rb���H���5��=UPlAm��PJ�J�FW��`�[���8Yp�[��;syW�ܛ2,�}�%��:L0�2A^���Ng
�9�j��,WW\,o=X@���X[[x,��B�J%���63�,�V�J�_d�<P����(���r8?P�|Oo�v�	
��ȉ�x�v����\b��ќ�?�ޚJ}nn�MAB����,��K?1��������`��9+�"ݝ
�ڔ�긭��Iɣ��	���}Q��y�kF)q{�FWZ$׺�ҵ.?�B���l >�F �פ/�c��p���l +9��hD�G�ɏ���u��kd�Yx1&��<���������a��x����~F�'NJZ1��N�1o�5���d�xCݧ�_�������H��b�����@��Ÿ�=�}m�D:�kPYj�r�Ucp�f�hhH4����+�w�q�[41����@.=/��|8�W����治7U�Y�G�^�|m����W�a�-:m���'E��t��f��7�w�.{G�������YRԓ1魡���4�~!�ف�� ��m�8,��n�uSDT0i���_|2���w�v�]]����`��^��$�8��W�𹡎�s����)�ց��&�]B�Q�)�E+����/��1�0�����3l���m<��r-����'�}��̚�)��ԋ{�h}��?ph�D:����M��(CB��?F�F�a+U�?*�ޓ���]����8,P/���_�hj��R���TL�ԏX8];L��X�Ѕ�G3
���A�\�M�=����̢��)Z+��e�@�7�)��I'>��.�8K0���<C<:->P�kTT_8Isp^4#vS�ش�e+�B���B�'ٷ�˓X�y���䌈0�7�H�FϔR��A)b��C�1�lŅ������
�Q���^m�@��Z�V�7�6���F���F�$��=EX�fU�|�?pqL"������R
�=G���h;��:�"���S��١/d��|����#<P�T�>��\"�4tmH8��H�K%�0*�����>	���h:�sR��þ~(,�w�KH(K=�bH-ǽ}�.�{3R�k�~n��
��☋���a[�Z+�����7$���Wlƀ9��PA���]�`FV�>��m/z'�5�3LTj�-de��aɠ��뢾1w��&��mN�Lk�R�ǪZ��N���������ŏP
����������ؒ+�4u�L�|M d�$���Y�x�O-��[c�)�U�M��œ>脹!�������t�Ι@�1���Q��'�$�?��^��U�v�7�帩��u� �m� ����DCF��\�Hs�����!~�_�+��)r����P�TQ���~Q�$&Z3����j��)���>�JO�-H
�/w}�}�
�X֛:��ϣ�-�]��:AG��dBO����z��ʆPE�Gh�/�H�dS�v�Pn�������pߓ-i���(*U�u0?G��ߥGpX���3�"	��|�/�5��9�� ø'ݲ�����Ia0�ώnq��'H�;5d&5{_**z!I��l�q��0�EI�� �|����=�#N-E
�V�g�T������[��T��)&��k��ٲ`�}���-
��{�dU;��Oa�A8�U��Vι��1s�������'�?͘���<��LW���I�+�&��i����u~35�mRw�ﾊ'��eQnTp�ǒ���=6�1z$��#��C��  6�ve�Te�m�"�?j�py��פ�1�!mt@��'�C�CW� H��u'�؏{��=�'�$���0��2G)�a�����r�|�	�+^ѧ�������B�%��,p�UJ�C�rh�Q�`PI+f������1�{m������$��_�
EI2��=,��Z�*SQ��p+QQlD���Fg�j�g7��ѐ�XM�.����Ӫ�ȃ󡍓(
�0]i�_��`����W[�j�6|1"�D�_�~����$�q�cU�փw �幤�,~�"V�T�w�3����M�%
?�I�D`	��vH��9�Y�h^tT���w���T.��E��~Qb�Y'\y\�b����L�yg�}-|����dP��'</���!���^g{��$��W%�ˤ�āue���F��e� !����O#!g���T�	���3:��0�פ���oO`�Qti��D8�l$}���Vh�n;THpN*!�5 �d�3Վ*| U����\��{ٰ����xb��(v5�̥cfS��4���D�f�{-�^��s����j��\��CBg��U+�Fa]
o�����hH����"�O.�5�u���l��|��̭�J��� -ms�L��끼������+<��(Y5D3b��6{3��i���?�wyM���>n}~�%JgP��"�O��s�]�\6$G6�Lb��\��=Yw*�*O�n�&�	]�^�� >�;g����x39y1`���4c�ۮ������A��?���O�JEc~�'�]̶�8�`��;� �#�&v7�Ώ��� @���"ʘҁLЛv��w�L@u�e�$��+)EU7�!G�R,�ȝ\ͭB�ֈ%�Kϋ@A�Ө#�b��{m80���p⒃Q ���v�w��P� ���5{s�>���~"9x�KQ���pgV��wN�7b��(�F?5����������|f��{�6S8OZ�X9x��w�Q���Y��`��f����y7$��Y>�C
I3;�]H~��	�\\��Ff�*R���P}��Vj��}��$�?5$D��
�9��]��K!��2��A
m'��]� z�����o��r����4o5g^2m�G���5����OE�E�EB$��y���'m��=f�����H��F��5��v�u��k?�7���6T�����b�s���m�9ЯAE`��7�������)�0:�X��ޘ>��`�ZӚ]ܡK��~�$�ۇ%+�?|Lj�K�"���e��7ڹ� ��W�I|�;�@�F�A�V��uD'
���*��Ju"����.D�qFX��Hd ����ʆM�z��e+s	A@^���3&JGfӥE����x�X8DDTM	,�B��9���n�yj��#ӃM�)��[���+���OyQ��N:p�T�Ɇ�0B�1��b-W��\k���b:�'��s{�H��T���d�Ka��/� ��7��� ����5�5������C�́yu��/�6 �z�Smٲ�;fן[�l��@ "�&<���E�~�U���4
=[9��l��|�����!�����A1sk�kl�}��[���9�c";q;���/��ݞ6��A+���eے�^��Bρ��;\��N�\�竵��;UV�y����|�SˠK�W�@S0gIf(gJ[��][�u+��Ӕi����D��E�	����(J�d `rG�?�Q)���&��<5E,�a���sQ����S�_�9:�gC�8�z�%ޢ� >N'lo��`�#-?
|���#��!�%U�Cc	N�-���4�S��6��K.�$��\�Vy�.����9:_�l��쌴m|a^\�t�c+�I@�:q?���#\�	��.�#������O�z0 9���"-�>)���bq���m����^s|G�~�6�O�8��Bњ����8����o H��~}��O洣�t�ܟPf��h��������tԚv~ڴB��p�i�ݑ--~eV*���V)���"D�[�8A.��t��������tF��ԧ�*�"�R���M$������q�ptB���ռ�(\^�B��,(�M�d�ܒ{x)��z�.O;-�j{91+��y::`ɩ�oK�I�:+G&0$�g�|���u�rM'p�̮�G�����a��0����C_��'n������#�O�|"3�ĕ��([�P�,����o`i#��
����ǌ�e.o#-Ç;s4��T�������l�b# �c��:�O�?���)��By�St����BD4�W��l�/�ktuym8�<]�3��HL>=Ӎ�z0�Y�"_ȩ�4,��e��Z#;y�>�Ǿ�v��P�I�D>�.��2�CO���3j"���9�$��y���4?a�9����@K���&3��~;3S�\�fQ({]�`��0l8\䖉�'�İ��z���A8_섑�qR#3LxLx�"����7����e�u�l��Q���)��"m���hsP8�c��(*�Bg���Z�r��K��1�o��U^��]\Ǣ�6;X������j�T�����W�E�!����}�	��]��&��Stp~j��r_�`݆z�̑VFG�0�~��v#�qx�-`�4��a�D|
��3C���ᄽ�!����&����@�_�se�r�t������簳"p_����k@	M࢞��n���K�9�&��Ø纹aV����E[���b�B��߅P��M����ٚ��q�X0� �$��̉�	B%$jV	���)Y���N'�1{�OV�;��X}�϶2��Z0�sO��] �a�!�x�^����W��M������y�B�s������,�#�����WZ�tV�4A���K��Zr=4�ZY{ᆟ�`/N�p���wvZ̕�8]�C��"B����P��ET&��+C�=KKQ�PX���`&���~���nc�m�+$X�r+�ټ}VB�AK�Xq@ciS�H(�|{C��W�ta8>����=,���
��1�5SҌdg}}��-�T�^go��Dy�*�\l|����i�l
�j� _�4˥�����M+�M��nq,ޖ��0YtP�;�R|��8atͷ�jwQa�L��u{�iD�YP���k��,��+������+tQ�-��%���7����B��1��l���*��1�Z�!hz�u�!��f!'��ybG���b`i����9t���A��׃=+D=B���i�Ĥ�NPg���$��ej_*��ɬ�.6#5�CZ�Y�<�?<�9��Os��Q�ff��{����|�,�W$b&�:�O���odF���d'�x�am���j\�)0%������$6����{�x�B��M��#	��衪 ��?�k����2�Y�!��=�uȧI�$?�;���s��6�<���]y e�M��|�Y�Qi_�?�%܌��+����(��q2�xn�r���e�0�6��E���&��5��_��ͬ�ί�"�Y@�s�M���)�����9F�U�Z,��,k�2e��?8�l"Wκ#���e�a �yy,���]��L��W�C����U�lxm�A�����lAn�Be5@@�1;�~��D�s�䨭�@e��@<�C��`�6U�����#~K��\�VC��O��&�k�j�ĽA��G�켘Z
Fk���d��n�Դ���u�t�ih��A	!���z6�&��R�D�k�"�7'��)YU��mr�����7ʵ��d��(B���OUٸ���S��Hh��|���xEw����u,��s���&c2�����J��n&.���s5�i5�{�X�ᴑ��:`�)�+�8�͗�0��w�J�:|�e�ʠ�0��I�ـy@I��вiCg��]!� ���~�<�n2�U�%�$��~Ýc@�
���A��l�T��E���XY�N$��$0m�XH���Ƃ�,,�f۰�G��yb�}�ΛpеlP���E���Ey�m��ċ`��"򶥝P���U�mB,A��>���L�bd]X"F̙�^�䷇�Y#��۾O$��?-����2�	a�Ձ5:.���PjHt~��t�!��Yv��u�5��c��ќ�m6`xW3��W`~���S�����Ø�\Q���$I0���B���ʚCk4*g8++�����D�vT�nl_��e���Hė��9Չ��_Y=�]���{nqn�#���_3���.Tk�w���`J:K����*9�Mt|�e&��x7ƃ`��O� ���Ƹr�a2	��Xa�Rq&H��;	�w� Ue��H�)���=B��).�J��9�	*������X{��\�V<�V�n��1`��%y�2;�d�£闗$�r)�q���,,Q�����h��3�7�\ؾ�!�&��9u� �=����Ь��8��zI�?A���h��s��ނX���!���~)��?�+��W��4x�!I�����~� yx����k�-1[~��5������ks���=5�mr��c%ad�8��٣�X5Izi�A�MMh1&q� |'��{�.�JxA� ��y=:N&�آ���8���f6�Q�����vD���7Y�"�0��L����B�i꼓�4Ү��IP����ʼ?�����t���tm ��}���N��#X�����Y#ec�P&�r)�Jc�8'��H���6������/~dvL�,c�Ǭ�<���R���C4"
�dl�[��vs����Ը_�֗>�Et�ڍjA<ѻ�q�PVbU'3�i���m�G���G�Nx/X&" ��1��#���l�~,U��T�Ұ�
hS9�FwJ�1��p��ݨ�G煂(�"*j�Ly�4q��&����ob���3��AԮB�GĻ�ں�3~�n���{I��)fjw��-ZP?�����x�i�Fz��yr�"kg{67�T�&4�||N^z��2���I�P�K�ͮ޼�j�T���G�B#�:p���q�;���]�����(��5��5�L���Zi�z�V��]
��zzX��;U����>O�SR�n��{��p�(�^fӎ�Wh��!�l�q��󋝊Np9��T��%�U���.�����=9�f}_�����#�xjKӆ=!�Αߵmiا���Cdsb2Oo	P)�s����;#�����u&�>.��.�S^�4"
}`���uk����i���p�._Թ�W�u��zw�8��v���vi��Ӑ�#Q5#�%��e	���|�|X\O������^|/�Μ����]ӟeq���c߫Y(�D��2�pV5L��9�>�~�n�i���<o$)ַl�>��g`5��~�~��u���9�u���悞T��ѐ:�b�Zw���-��&�Y���Z�4+�F{����LyZ��ř����>fW2R+�f/Mn�b�β�RYA~��hR��AҪ�&��8�B#��]d
�h2\�;*ߧ���N������#�߾M��x`�[	P�p$�?|_*g�``:�UZ��W�th�|I
��ٓgtYת"h�-K�a]W.���ퟒ/���?t��N�������ǧm���;H�{��l�0�k1��{�#���F �嶁8\w���4 A�aϞ ���s�c�j*��g��Pf���+��a�<���q�B���h�Ȱ�pUH�/�ńg�hm:,���E5^#0��ث�v� ���Ҟx��ʹI��} ���8����zi����e9�*p;��(��P Bi�^��Ԅʌ��Yc��?{��ɇ�c�c���j�}���q712�SH�����R�����]Y�J�*��ཹ��������������}�
�l��{͆��,<��+�(���&�m=��I�4�����!�ʠT�S�	�V�~�S����;��2h�:��z���`�kj��}qߒus��)�9��(x_��w:x���,��?x��z�Ⱥ���p>�B�.�@-�I͓hQ&*�����Yj�뎴5���*7��ʎ�Mc��&������5�xp��8@�/�e�{��/��gyYDْ���Ԝ�}��������"M���	��21T��3�dS�}m�������ht����Aʰ�[��L�V]�X��]q"�������0�_(}V������7/&c�B�gJJ�ϟ��I���C��U�I��@���O��vnpD��)Ԑ�'���[}�e��ׅRV6aa$���qmtB���(l�?���`&�I���J�v++���jO>���J^V�c�ͩ5|��2!�H�XG5l��:1�@��.����q�<��d��#YI=WtM�\��G�D�3��^2��Q�kH���¸�k[��ogh+ZW�Š��:�B�iqQ3J�QN99'ue6k��	-Eݍr�Ï��)� �F�5�t��`�޽�� �]��2��	5�-��y>֖� ����1�!1����Յ��0���c-���{�M�� S��ֻ����A��=�� ���<}��.e�	}���	�DV�Ձh�� 6���s�5%f�C�����#(��!�Ƃ-�C!��g�d�?�~uTS�����Y���=�?r�b6Y*�n*��w
mη�̳�4�{�#2�ִ�P8��E2���fZ�w��NN�>�LZnJ[{/��?��M�]V��`� X��1�n�5����R��iV?�ؑ�հ��N-�Q��C�/��6'�A�>��O��3d���/�=C�#�FX�t�}��JP�┎zF\R\��8o"��p<���{���R�� �+������5O�ϑ�y�h�g4��jS�NQ��^��OrI��zO=��»a�1c���������©!gAf��؃
`�,�l��E�&$|l��<���Ҵ���2�YR<�
j1b����g&�<����a�C���t�E<�,�\�I/[� �46��9^[Y�!��>��碋�@��.B#�ݦ?�[����r%�+IFV����8t����ѱ�������8h�nZ9k�23��|i�拌�oh�$��. )�2ъe����v�b���[���x3�|0�%������]���5���1��`5V� sm��⋇V�nP����3��i@�Q���$�G�<sf�el|��PE��7�	�tD���z!�`@��Cp��PH(��,�wQ.2��#(��Z��I�V#H�ea�hv.���u���[�^OU'E�=t	�,�h�=f1f�Q�Lj�~�f]���>�'�CA�
�MA�2}����Nhm�2i�N^@x���ʣ���^!T�e���2����E
�����<���I<voN�K�H���N���Oc�#J�#�8&܋���'R�0v�á�/ٴi�L1;S��[�����*K���S� t,|Ը�P�ť�X-l��6��W�k��v(=��KT �47#�@}�h)Z��`�b�:j���*J��{�Y�{k�?���٠���4��y��Y�b�
Q£�~t���s��Ї��9?�b=z)�<��f��d�-
$�J*y: <�g�jss�!ې����E��É�%W���6��l8���ڨ)aZ��-�Q�kT(-,���;t{�P_����)/�V��"@/�f<2���ɕ���t����MQ��i,�ɚ�� �f`��������އ|'��WAU��+d��gr�,�Ezg�*��G,��WUJ��z���4����9��?�p�(���ֽ���0�I��lPTɬ�=>�4M����fv>q0�y�U#	�����51[@Ȕ`a��	�D@1�J��������ϵ��;�M��6��W�.Ζt������ ��Ka�T��$ ��ΫF-5m�p�G�3����R��_l�����ޖtU�v��������e�Ǥ��~W�<��8���#"��
�?�3�ɏ��&�R`�gDޙѳ����,�&��SW�a�4��Z|ʦ����)��Y�z��fj�7�m���Hy��ϡ������1���Ag	�i`9N������CC�/&W��`E�:�OG�6/_���æ�gi1y*���ن�r�>y\U�#.�C�}��K^aβlh�[ �%�9��L��\�9U��q�����#�E|��>D�Z��r�X~���ɠ�I�m�r`����ϋ`�J\���+K��?��[ʯ��4r<�D���vAE|�(��|�.�ŕ�������BI�k,k� �r^�����a�}�ߩxfy��^���MݭN�R���"y�7@�N�����:k����nS�D�KH��S���:�}��4 �q�:�9c�ZZy,����Bk]�k奵'o��g��yퟟ`���	i���~E&C���V���`��?"7JשQ5�ܞ�I�� 5?ޞs�����$�[V�bIG�?�.�l�8�&슡�b�Ӱax�$�*T�=�5�\���g&;F	hZMQ'�����J��q��x$,���~�3�5[!����y'�f2�{:���w�2/�
�T�4*(�P��nae���Rk!bJ[哘�b�m���s��@'��T����ˇ�T�Vo/ui�ѳ!4��e�C�� ��tn4`�d����N���:;�����^T�\��l�P����J{^�C͍l?-���$ډ~�	#ݵ��������� U���]��ɛ�(|*T���mߥ�'C���*����m�Վy��ܒ������ou�._����Զ'M��,mh�Іo��/�Ĝ�%� ��/<L)�����(�J�)_�]E��pHC�26u:粍��j�+A&X��\�E���y�, OM�Mԛ�8��O)x�Yz8��y!GxR��x��]䙯�6K���~�`��^?;��4��{*,,x)�		ɹ�;_��|��d�Qv&�7��\��a���O��r���.�b��w�4�!L���Ϯכ�3�~a��ѩC���S�H�{-���vdh�gu�a��"��8������*���{?��Z�)!f1+/�:}�?�������������m�0хԚu��j?Ou���;O�>b��z�#��eYa�Q��!0<�Os������#���M����ۙ�J3J�`>�&�������.|� Ʈ�eP��њ;��c��G)��H��%q�:�a�ĦpGz��<��z9�PN"��Uv�5~��Ɯ��{"���sZ�;K��ɤ�*�a$I��!4��̢G0�,���)Ms����?g4#�����\��Lw@ke{�5��i����L^�P��1��JWLt�V��j �kI�a*%�q�l���L�SlpsAB�/���QDQ��4$Ϥ^Z�B�r��lHA��C{������ؾylm������S^iz�s��v�ӑ?3.V(|P���p0���q��F��N��R��ɠ��w�7Li�K=k��F��;�rF�T&���\$|�>�ω�%|�h�ʗ�CJ�cTx����H�6왚�" �6rb�t<���RQyY�� Ӷ���Á�)�̔�P��m���6J�6�P(��bp��>;Z^3M�I,[\`����s�&�Q�T����.��>H|�/7�
�w����j*X�����R꧵���Mހ�U�!��63�Q���t�X��w�[\���G�ZSv,d,�\�����ӕ�N���LN^�<m ��,�h��t�����ߗ��Sp�z'3��^�j��ٱ9�9\9�%鹟+���&趝D�m@}Y�����K}¢H�x�:����Y��_�\`�B%�upB�n�u��#x̵-wmQ�1k�T�T_D�ԛ�^w;G��[`��`ژS�/y�-s6�ǎ"j%��}O�G�߮s'*�� �Ti���HmU��БMU�AEG�ޮ�mا���9����|	�a�����Y]���^���3nzS#��'���"�̦��e�U!e7DG[0?��9�u��3�_'�C�lt�t�:�Cc�[0@����k�>�b�M	���s�͍I���ʞš�N EN脻�
�D���2�����T<�N�K�7��%�#V���K�eA1��1|�n$d�qؖ�b='��}�UP�Xb���^t\��x�W� :t�+!��Ħ3Y��op��8�X|gN�2��h�;��XY�XA��/�B�]��Q'��в�E����v�ϿE�Ѩ<�ASE�p�±����P{)�	���2T0�p�dp9eU�2w��▥�=��X�R8l�#]�B�Eq�ff��ʉ��p<�\�;H"Ȱ�K��m��I���d�����m��-�2�~n�"r�ha�K1
=��T^K���{���$滰�:5�2d��M0� ]�ɳ�����س���#�1E�Y�n�� C�=A���u��_4��s1t��l�ܴ��2���}�o��H�SȾ�([�H=�cfT�S���W+�7�0����T�0�}b��K��9��:��pM�M�g�}L�I	��(Ȩ\�ތ���,N��U����/)�yFq:\��x�՗r���[�|P�� ��Ѝܐ�"�2F���%<�	�e=���خ����K �Ϥ缱;����'�U�(��Ŕ���Y���Du���Q~M�`��>l����!�1
0�D�y��%^��M���'(�%�ĈL��|1�q��J��:���.�%~y�ǽWA�<E084�v�n��־&�g���C�Y���v�O����R_29r�&(��E�~�$B�KR�NpV@�W>ka�<�ߜ8������P�^ �[���d;̝��K� ���CD&��t�3<���o*�굹H��^�@(| U�iC�	a0�>#�hx���pD���y,��_Me^���R���J_ZUh>���G����Q���	#�hz��y�!��Dc1�������t9<��������_񺪃4v���?�_vؘ��Ԛ�p��+Uƒ�
�<R�2{+�-���}��ޟ;��p��f�㯝���-0�7�F�{�8�K�a!,����ݥ�����r��RV�K���6�.惉;�&z�EPh���"H�������}������(5&Xls�|���Kyx��4�C|y��m������cw��rB�A0����Лg�N\��KH�x����ۗ ��+&�0��@T �d�	�:ݹ�������Q��w9��4!�)���{^�vO�d	[5t����?�`w��#���E'�� ��;�Ԙu��G��A�ί��+��Ͱ_eP:��|M��6V��"�>��M�		��^ߵ�~Jot�5��߸�12��˛��߁���P�)�<�:h�H����ٖ���:��,k��$ק����h*����'�N�?��е3+e���ċ�
��
�Lf�K����P%[eV-z-gS��Y��Cg�K� �*����ߢNO�nLT�;ML6E�zЏ!~[6@z��͟S��{��@��G#B������F(�r,�X`�l��䚶���q_Ʀ5��YK��8��^z���'������4�����>�������AC��T��2����K��u�� h(L�Ҭp��	W���S�����zޖ-��L"�#�C��f�nI���+9�oo���<	ӻ��*�!i΋` q��~`Tݶ_P�J�Y����ƷAM1�>G}�egYC��bۀ�Ĺ;p��MmE�ӹ���F>�u��x�Q���������ǁ�כY�i��d��x�2�n��O��O#�ܞ	���wUX9�ݴb�n<%��oM�\��0�D�m��2z-1������NL��B���o���A��Q��ť)<�@��M�r���xZ�:�
o�>�ūW����l�f7h���|��FR3��a{4��vx�'��"UIx��7~O��B��'<ƺ��:kH*����%��e=V(hϐ�[i|x�n��YaBdi��ܳݙ��Hh��&�P=l��y�AQt��k�_��5��=�L=�h�*Y��`��֐��Ș����%��0A�-|Q�p>�a���g�#}'=A���ROtps������ъ`J�R*|gb�B�c�f�$M�hk�⎮֯����95$��u�6@M�[gg�x�`X��~ȵ���J��1�K���.-�#��RΌg���Y��!�ABlߋ��XY���l���s(2�錷V��kp�(?0�w�񯳔��DN���bT�k�@s)��O�ٗ��O�>��o터��z1���A����[��r��i�DP��xʷ�Ӆ:��d��]�g�<1;�k�(�P�0�0+�}��T<�fY1����4�W7u��n+&Okݞl>�8CпT�
�!�s�@��8@������̪�U�|h���!4��+`��}rqz�{�R;�2�"��χ}�ַ��F�h �3�/��F(si/�J:�0�3�5�mUm3��*�s*Ȗ���8 �S�f�28��0�;�_�~���B�,��W��=�J3j�Pt
���_���`F;{��O܂t��o�NԮ2��s$����<1��$��*Q�ƢN������Ɨ�\�	�`�I�� A�z�!�6��J:@��8 x衁�uV��
��vk>���RuW'��Re���2&��ތd�}Z��
��M��ů}�d���>m�B��@������ZQ	��?K�sR������@<;e��x��	���1��m�?~Z�4,#�����z���
)=#K	[��t�8�8b��}zʋ�i��c`>>ZT����d� %iX+���kť�=7��G���R~gp�YLgr�+F��׬xi�6ޫ� ��oS&���hB\ie�")�_* �>��0H]Ϋ�}o���� �	��E9[c�T������/ݳ�}LR�>Z������<< ��Ʉ�]�t)	�N���_���� ����̍�S�E1�>"�a��a㯕v�ۊ�h$IFVӠ_��P�K �V��ɛD��mq��2��n�H?֟f2����=����@,���lv�#pO�����k��s&Q�%��.�4<i%�{Yf��O��ߋy��ĨY$������rR��'wZ�����27�]�) �ff����0ֻ/ ��'o�-��;�O�3��5p�빏hLS�N��i�ꇿ�Y^*c^� ���0fO��].�Ѣ�='֦@��1O��ЎR�Fl'���E^�Rd�v1���N�J��m���^� '�\�)�J�c�:.#��5�hu�|�$	mTC ���G~z�9}������tO3~�V���K$C��e�q"E�8I|����5L,�j�C4?%�[�V���m�U�;�<����n���u��i;;N��t��kx�m�E����d[�-��<�Sg[�F6��&	J�п��w�Lŗ��x�Hգ���S����=���j����"��,i�ԭe��5�pg� �0�#�˸V!�C,.�������:���\D��l=34�������o4[5>;"�#4TC��2��q�x9K/���Y8'tR��k�(:JP��,<:��ex�C�v�Z�P��u�[�*~La����	��K|LT?���H&e?}�!�a�8�/m
@{'S��*F�U�+}�v΁�]��;&^E4�8L]�ôay�>��8&�b�#r��х@�6}%��>x<m�+�����|g�����rx~�x���E��]y4��y�������0�$�}\4hp�!C���⦤�:�ׯmXu��Y��,&�����8mj9������1���Y�T�to"��@؊�;���������<��q�ӝGO���z)*K{��"��%ӡt���Ւ�T�vd���1q�k��ġz@X.����,v}j�ݥ�{.��G���n�ʳIƯ��m�%�é��Y�V�iOV��y��%j��g���K�Z4D7��93/J�^*��H-m�V
!'�j�_2�j}��m���)йO��̨M���5V�щ�?���9ӄ���%_��w%a���6�T�ĞC�{	��������}���'�P� ���Ă��a������S�U(R�"P8�g��KZ��ؘ+�]�x�8�<��q���%k�j?g_�Z��ABB�]������X�9s�	!Yw����S�b���¯Qz�l�1��~�w@n�U���oPk�l*��_�z��va�D�Nu��B.���,@=Y�J����5S._��剹~���̽KK�����������/b��5��r*kzXGim��b�X���%��.�3y���2��oǶ�	:/���oRd��H{�E.�mDb!6Ҽ��{�Z�#O���矸����s�-D���Od�0���J���󶎳��2���z��_�����S�n�'��|��淙ٓ��56k�_@Om��P�?{��+�H�&),~�c]����&[#�6J�]bF75@P���a�5�W����=أ���)"���q��gF���ѕ�q;0���Y��U��	"pwec�}>6˛����I�P��RaQL�D�]���']�l�B9\/���ϝ�g�"M�\�R�o$���~��a���=��}�@80}{�B��|��oP�D�Ik���������Kbk~�J����1_qy�q�͋�`���lh���[����9����u��+ݏ��k0k$��K��Ȕ�ba�d�FWq]�%�X�r�
h�7zF
����J�e���tg��*DJ��{�?��"A�w��,��j�P�كY�E08�#��B�t�������,
��]��M3��i޷+�]�օ�ᔼam1}^�Vʕr�x*���DB��Y�hc�G��֗ z�W��-�gEu'���/�v(�HC(Y ��1T��At�6�T�t�`��M#�6:���ILI���	��$�	<Oǈ��(�<	�|f��+)�X��ʽ�{2tt�E��s�H��gE&����(W��R"�>!^�`F��h��r���,�3��D��Y�A�,4B�Y����f�m.�]��'�ƀ���Ukbw�m��z!���wo8�~��	k���āƽ�TT���5�貜T���r���d%gj�.N��Ў�خ ۝:`�6�^�j��ch��@p�"g�Vֵ5|�B(R�tԍ�7��<��d�!tFa�FH"V�!(f[_�\����/�'� (�;����s�j|?कi���,�l���{�E"��ǰ��c,��0�I/_{XfJXU���F�b��|��6r2�������H�b�ZYV���u����6��>����h����=+R2�8�',52��Qt�or�Ύ���
����?@"<lk�;��0�m�����&��פ��� t^9�_xi��I¤0��a�V�b�f�d�Hm혜���&�������M+)�0T7�v"S�vp��ל�8�FO�q��d�m�F�Ԁ� �a�p�Ck��:}ɇu��n;�����Jqm��ӡ�Ee�$�,�i�3kt�����jW�R�e�-�
��bh��p��F�Ժ3Lc���Oz���iX��a�=J8��)?�-����~A�>i����gS a�bhV�`eik�>�6~�G�>��l*D8��i��I0�Uk�,�`!P]ą�n>�߮�?�P�T9th;��8��_WH=��|
C$�]"F�=O;U�-�,i�������
���c��p\Y~9��1���*L5�]c�՛������%�" � �)���)��_Z�SQ=�x��-��B�S]�{N܁M+tܘ1z)�H~����J�-�۠�&z�a>Dr�Ch6���Hj��	����|'b%9�:ZÛ�˼.���8*�k�� Eֲ��\(�B̴Rc
��2hx�D��'�څ=�OQ�q52b��8K�*���"Yw��<,��hYF���/~�xc��P_>���)�q���k��/߻f�+vt]�F��<`/Q&JFVׁc���4[]��������s�ʷ�j�-�uv���I�_�G�����'�vμ1�i���r�����+�>�zSȧ͹�G����0�cT�(����+CS�J_�{@���A�?hu	�ݯ�(ӂ�blm����,�8 ;9�VNN��[���z�� �F#��{;+s�o��=��s=�n��}��q�A�a�3Zȧ��J�8����ˍ��"S����#Ɍoy3΅��Gb]v�rP��,��l�dr��g�y�be�hj~���_�[ϧ�}@k��e2dČ���4d�hܫ�[��I�W�cQ��Q�ኚX�U6�i3�m&�֛�į�P����r����`mBbKb��ԯ�o�ט�c-VK�1W?���$���p��@e�\O��u���OdE������ld$���y��>���*��\�صhQ����$4���N�2�SȌh�=����CU��q�mn�S�|i�u /t6k��t7@/ �[��	5��Q�Q�5���}
%*,��*�F��1ۇ��!q�P}�,(S=b���V�^6}X}��42�l@l~��{ڬ3T{��#��Q��dd���xi��B��ޜ�4��EPom�c/��1�;�j��fT8B�����U�!;C���*fI��`��u�]��;������˵%_����Ý�ͽM���1�	��u���+I��/���u�D�pwV9CW�(VB�aN�nP���tp!\�o?�4Q
 kĎ��!����D��ί�'!3fJ��Ҽ�}OH��M��$�-Xm[��.�|9ՀPG�[�;*�I$��ܗ1m�B��:'��9���ϖ%P
���TZ��W�q�\��S`F.4��� ��i}i
�ϔ�/fJ�V����f�<d�>簬����=�R��~K�AyB<�d,|`�����Pt�}ɃVW��|g6��p ��:n�����1��g���C7�_{;!RU��o%<�mo00�C������;�=6 %/JXc���	O�1F����oIG�Ye2?�b�B�^e��:������V��KѪ��6>��)���]C%ፀՆ��3\�a~/ZK���Ԫ�7���<@���~�9�b�@�#`|� !�Mc:��*+$�����HF������O�U��Z�/�f<A����0��Q�k�k�6`FN�D��J�{w}х0�&"Mն��Y��$�gz�d�и^�^Q��5�+�QǔddKK~��R���r&/�$!t�:�Z����$a�=HO��U�k5l�\7:�-�F������π�����y�e��
�o=�j9�[=��ߏZ�������3@dq`�����DN8�
7~m%���.���'����n'����:j�m���s��p��͍��i�@�Z�N��r�b�+0��4��E����(Q�"Xm��z}��Qg;���J,E'��8|�g�QcN�V5wCdT�e4&ZY66�O$c���HZI0j�5���_fΚq�	m'�M�ۍTF��@k����f��?�S�|�争t�u
+��wĦ��.M,���2he�X�k�~>ZVq����7�:����*�餞�(j/]�{�G������N����J��3$�4���ꅲ��k�#�*��p�YY��p[j���r=�I��ܙ��5��C�]�ZմITz܋�N50���W�#[���[+�Zi3i���2���Ո������X�K�v�},�����2���U���d��y�4xu-/�H�]��:ǿZX�p^[�Q��`O�lm��(���6����I��;�3�N���իtk>|����,���!��|\�M���G,US�bm���������څ~FҎ`r�w���!�;�c8�h�$+~�xٓJm
f��su� C���C��e�R�!�j�s'v�x����B.�߁s1lz�^� ��o����Nu���k���cF��w{���b5��}=FY5�e��Q4��s}r�?ʷE�}8e���e�-��T�2ґ�ܪ(yTR0�1��]auh�^�އ%"˟��'�<�M��2�6�5X.���o:�9p<Ҩ>��D�#)�|2��ͩD�l�
��C���2�:==�}�bFe�Ԉ{�������c�=71�WcP�ls|�L�O���gͬ)W�})�S�^� 66���5�E�0B�U���,��ot�=!���e���o�b��^��5DUAw��P=^�w��ꠂ�P��rI%�k̖�/�� �m���a4��{�]Mn��v.i���}��G<IH�6�R8>\,M
����$�ߖ�_�O��-��T ���\Iz��#�ț�6��t��N�����3�@�/���ō�5;('�0�䆂R+q�D��!;�U��EvG
�Yh-[�Mu�ku�6�ntb�p��́���3)����2�3܂J_74�Q��ޢ���������	Φ�Ns�>-����H;�hJh�Y��/R<A!�����W������9y�)Ӥn��80��9�Y\�(v�o�mm�9χ+,��M	@�_����|h����V"<ǆ�L��W��#��8�X���tjhGl��t*9Pr{���F���`ME���
M�D/Ө,_����Vw������E�{�cZ�o�9s�6�gK�pi:�� k�U�;*+���I�gr�ș=����|$.M�C�Z��VU���C%'���k܀ϏnO�@�tl�F�D���Λ)z},l\Ә5��L�D��Sn��A��� �����Fδ �G('�=5�]��e���7G�zk���I$T�삇"k܏_|Sw�g�  r�r;�c����s��l&L��0y�d�30�昨�"4w�7������N��W�y,�X��nWy@�)�N���!	w/И1*X��y�oME�r�a#~#�G;ol<��C
x�l�j-3���)T/V9��S��FZߐYq=�
�ˑ���3X3B���ϸw��Q�(�AYO\�.,G`��9nէ�L3�h�:A��z�zϝ`��R��s�����7�b�l¥��f�*\�鮜N�ת9lX�8��Z=�F�X�����6,:���r����-B�QˈOT�l��m���ȿ�xx���Α1��m��T\�36L򕒭�� �B�	�"�4��f.����f�Y��������3]��eo� Z{/fT�Y�ػ����͙OV�1����g�Za�Aa	m>l�m��x��+��6]��L;�բB茶�s���k�~r�
�����ޭu��ң���'�3��%k}M�ݮG�����G��&o!&�t�A�gP2+�"�i�3m�E�����&�����e=�uz�@1e���z>�ϲ�ŦE-N�V�B2w���,��P(��l�FL�g�p�;��7p�b۳�E�씟r}E0w䑷JU'rkM �4�A�\������:qr�*Z������]�9�)2m�)�枻�.�x(:�q��f�F\��NQ�FY
�_LM���d�ة���O[�cş=)m�=���+��ϰ����r�E솞e)��ezJ2��`?�5�
}�]�����Ѡ;l�/#ώbv�&�f7���Y���4�WOLj}w��X쐑QU_��=�T�t����/~�}���"sV7m��fZI~`q�>ɬ����7�ҝ�y7��M��0����S�5�̰!����Y�}孊�U�rM������8ETA	��</��J��(.Y���wh�z&j��Ti6�xߢ1�G��t��ѱ+6�ln�k#x�6v��5���E����GŢ�fBH�:s�Uy��o�M>7��ao
��Sq����NJ��V��(����6h���"$�f��`��c�k��e�n�`(5�!zS�
�t}Q�c���i!�,&{�r�������߫������?mI�1!�y0�I4<����Mdgy���oI	�2�Vg�i_�:�OZ��d��S.�9u�`6�զ;�Wl�����٨�~-C1�
[�+��Ɇ��N�wy\�xw�{ v�����ݪ&W�ɹ
�*�4e�'���˽,A�y�D�k\!��ZgG�r�lQS���n��(�U;W_�a���|}��	���rJ�t��9����j�F�����U��Z�3�%V�#>���~J�<R��!��S��u��ƽ9����a|A���ǋ�Sa��֌�PS  ��hk�iy�Ŧ@����Y7Y�9`�?{j cEf�b�ϓ0�]�sTD�Rx��-s���u�'�[t	��ѩ{N�]@x��<����NG��e˸�$&�hf�C�	��>
-���yO��� @�Knw�&���~'�Zح�!��A�!�Y&<�rd9�z	�yw�5_EɌL9���S��t�D�p�NkH���Ѽ��-H�x�Y�����Ѫ ��w���A�֞��H-YN[��`�4�ܕX �=,�����v,�=���j
����u���a���/�VA����(*�ɫV�t�(:�E�G0YI��7�N߸.k�c�@��­���="L#�����ɫ�%����y���I�#����=�aѬ��~�e[���{a���h�s��	Y�:X�1�~�:���a�x*�����8��~��/�7N+�"p6)��-��=Ƨcm5�حV��	�J����R;�b��45pη͖�4/<!y�x�Dj���#�ҽ�[��iVp6��`�R�J����M�������k�dY���L�pq���>r}�{G)B�5/��V�7��'�c٭�P1�nm!:�\�|l�x���y�[D�)�-1R��ʽ���#8�?;Z��¥�|ܢ�m�����2tI,3B�*�����'Ղ��3B�h[������c�S��$N 朞�с!��J^�E�Q������|q$�V��@�G�}I��� "I�h%��*�ќ܌tle@Ѐ`!��a��_���}rt��%Y����7@Z�j���{1�/0����@s���[�ਐJe���U����0���:�פ�V��C�Y��sp�i$%����W�gx����!p�����-��j,��K
��?�����w� �cSـ��L)��jq��#_0� �����Nz(y2������Y��!�L���e��܎�v�#�@(���s%�M�P� �I���z����_��1ZG]�4i���0K���*��g`ݝ����]�����R'w�s]R�5��ʠ,C�4+�x�s�w��%ĺTQ�ke�c�k�>P=�y�G�L���p��Hh5�풕�d�AEv��d]��	�������傆��C�f���z��Bghu��]ĝ3{t���s�ΆJ���֢��Q88�;�
��r(t=�j)���[�����tYwi&��؎5�����rAJ�.��2d��B���[����Ǚ㊺�����֣N�CKF�7�$�����=�Q�^g4�d���������F@���_����C�2�Q�>�瘰�H=�
g9 t�&0o���C���{���R�p��P�i���C���1Y����|�8q�g������{RSR���e(�m��ņ���ɓ7d���r�V�� �ݕq.�B�9O�y<�@@�;�Dx��A��}��dJ�K�H?����!eᮁ�P�}{P#�
��n6t�Vln�8HjP�Q�;[Dxl�J7���J�@U���>ٚ*wh%<q�6�n��k{�ڠ^�/�
p���?5�S'5	��w��]n�A�r�!�؄���U �|�iM!\0L���<FG���Yr�Ӌ����b��~bO�hѨopW<�T�Ƹ���&Lv�4␷//�N�MWk��J�Cp. �
�&(=^�09щ��0�`�ar6����� ��*OP�+���6tÌ��Ub�	?	)����706���i��?�4��a�~C�Y�.�-��~�&_օ�� �$���'|���m:3�i�?c�ژS�i�ոT:�l�.V�J�#1��۰�*H'�`�d�Ͱ�mX��E�|�ݙ��G��p���0e6�ް�>��cW/bE���Iha��*���3�N�؋@'R���l���@�2��r*�9c&��0�.�����,�N̜1�Xi�V3U�&���E�,�����.�k��T�W���K�a��z�R��_�����+��3���@x�( ��xT+��x�����..o���Ô�t���R$-n���J�Sjzo�x��;n4�f{Q�a��3��p��?%��K&�5o`-�å��X�WX�Kb�C�w��!�N">�`��9`W:��UL?�Hڷ��W��|y8h���x�l��"}�rܶ���Z���\�`b��5-M]m�Ґ^�jY�/��F����H
#�l��٦�M? ���ͯ�e�<�Fn���up)D�-O�u���Y�)^0c����+�;@c�h3�YX���U�e33<�{lay��kd��"$�$@0BN@�aY� Z�:�8��b�(V�*w.	�Չ���v��"�u2�	h(��5��1��K?����rd�=C^^��rڤ�1��|�{��B���c��dL��U$� �_��K�jp�:I�N�`B�f���t}
��Sk��)�9��;L��0�ƼN*!�d��H�Ө�<�1o>F�I�A~ӥwҢoȳ��p�����!�˝�X���R2`�&`I��P�;��-w�	�σ�Ji��+�J��ysv�M�>�`$���U`?�����m����Ws�9[����/_�Y�|#�u}¿���_�u�,i)�94!���ᜱ>�?�v�g1��?�Mk�O������1�X�+���{S!�d����o��j0M;?C��W�Y���ܽN�j�n��e`�ф6�U�٪�V��oہ?��5�\H�m�##� x���ٰ?��3nw��z���7����ݔ��Djl|��)~��u�����:M�َ{���`�Ol���~��������%���>�C��,Z~�,���&��B[6�W��;,_73L�4^\�XTƆ�s��£�w�6�����p���B���@[�d���m3�+Ŝ}!�1�|z�dz���V�܏y(�|h-lM'<!4	�����*9�k~Q�P�$�hֺ�SU؄Y�b(�_^���@��\^�F��6�����(i�G)yN��[��329�-$V2��ۥ |��鲔�+�v�2��GV�)oq�"ka��Æ|$\�%���8E��2r��G�ԃJV��4�q�����/i�^Ή3tsM#�K�f��mqz��B�]:�'vJ�,�We�%� P����!��K��rhQg�dNL���W�I��y�I.#�����a��V�F#K���s=i ��uVh7�yݣ�۷S$.�TFo�L]��|{�rBa.�W�'u�[-���!�an��V4|ݷqU�H8�w���:K0.����0��%́'���_�+8�b���W�
�'��+�� �w�]˔)�X��=�7^�D�@��Ъ�	�Mq-���B�=�*�PI|1#�#�r�V�����D/"�Q�,�!g&���Y��*g�9�>p:R��6���,���O]�8
~h���e�m8:���Ţ����8�T�u!u��P��P�Nf��g��B#���}�t�
@�QSc7?[�g8�KY�4�������Ѿ	�䆜D�#I�J��x��~���:��T�_j#�, �lP����h���,��:���I�e` �����+���'u���I���:�
�/���8��F�r��`��x��X�v�>����ԌJZ�$�v�V��^(-�;������HеQ-ٯ6`C%�ݮv,��Gh0��h��`҃t�<��T{�<��iq{V$���)Ij6��~����.��#��a�\/g:%,���7��[)���`����q�'��D�R��/�`ȧ��t ���ք�
kJ���\�?���GM�2�lܽUoh��}Ca���z-�@���|�J��|��%���`��'ܒ	��O�Hh%
b�Q�TK�GQ������bs�����;�'9�YT���q�7AV ��:&we�OL�U0���d2�H�Zy���Ic�'Ď9d'~)y-1C�^!��R= �Z1� ��ӷ ,%�6K�^T$X�@=�a!c���m�`��}�l��9%Ç�����ΕY��܅�H���]����f����7
�sT͏���f�Uٺ X�S���Yqp��l2OfƏ&�3C���9���:����&0�y���e  �A���`�	���bH|IV��2�܀pL�����i���!5,��s� Rd�u�	b��=�W�KXS��F�-v�a��u�:��5k��"���g��6�Y���`���Y��2���	`B��dD��X-]�j	N�
�>�D=��+ENw�Hy��3�e�V��� �9���/t��C�S���fJ��9���f��Z^��o+\e�e�7KA<13Rm�����4|Y���q2�@�֌��g�v14N��ʁWl������?�3S!b:�U�ΩV�G�BXd�����3��]�-�nl�A/�ߏ��gا��v:����4[�J�n�O�}qs��8���`��Q����M$�굫���eقbk�����t<���a��vmh%�&T*2��Nf�x�,��){���BcO����5�����Wgd� '־j�LB�@m�W�u�?G��P]T�}^3�1�|G`�����l�HF�$\a6�%WI��O�JG,�޼-WJ	]H8�v)�-/
�@i��v��,��O�ݿ{�����Rl��
���q
Sg��
���hrnԂ;�-䳷�X�7gUV��)�~u?�Q�z�[����A'9,Y2}�[R�o�sG���ڤ����٥�+H!}jn=�ZnZdc�|��3�"�ǋs&�'�1���Q�S��IlVJüU7��<��4{����`���*,ʸ�!q"I8bXE1��5CX�� 2� .�^�ȅoˇEm�vv�9����85��#�!�p�,��'{�cQ���5�ɋ�E�w;3�M%����R�:��6Gm8.��.a lJ)$��zm>�<>����� 3�=�����g��~l1i�~�
���7g��ioe��tp)�C��~������ҁ<g���H�M5�?%��]\���j�;�� �)��y�;S�q���E>j)�:+~�U	b�K-�W���9�i����ޒ�tE��$V��f�<���)�4=�K���u9֔�'3��{��U��h�Rjg9���cҡ���g�UIR�#1y2 �ns���<�O�ps�%��Y7���DkD�P�R��ʽ������"��S�R�H����]�CۓA�1g��BS6d�~!"Ai��ۙ�$�Կӭ�n>���W���@��(\�}������-d�F�Ng������ ���/q�`V��ء�<�!�a�������2.���m��g�a�E������t��ͳgIF��ҥ�k�a����r[W��4;�}�D��T$¿�6H�hZ��m		a���������4�e���A����˯D�m/�*-��l�<��^%�^c�!i���A{�s��;���\	�]�C�ԑ��՞v�kx�cɀ�Ym��� �>r(����V���r�� t�_�	c�ة�)o��5��6v�u�,�U)�(�kS�|��x�<��_V����hIx� 2�!Z�Ǟj`F��F�ʳ�%�h���E�Uo���;��D���-��/\t/{�v�A��4(b���`��"J�O>�Vk�$���N|�����-o*nj��)�_����K�ms9X��>�Ǒ���2M$�._��&)<)�E(=��/s�gD����_	���,�?'N��o	D��Xj��k1�(���gpV���Ԣ��n:T�ΕS�@Yց�"�=��⤟BY>@�+�������7cCڕv�`Au~
�{�0��#���u���.R���K8J��B1��b�fPo�P�"��Z vF�U�Gw���u�����g�E*��U$�M�%3+���M����؀��nV�~\���G(���E���� e��P���νem'D
����z�oL�=�y��jOX�8�Ð�V��[��L��]Q��ʝ����é�����HW�� q��	�x�i�*rVtg��f��E�N�"Y!zm5��6��:��#��׹��������Ka����P�Q��%U�s§��R(H�v�3��51��c)[�[�χa'>�g�N�?I�;�7�N�_ȡ��h4�ܦ�4r�{7u���3��QϹ���
JT��jn�����#�͝��c������o���|��� ��r��ABp�E��7�|S��x�Jia��:�X�y�=8���'��e[��À^��pFQ�V�b����no����/�����٠pqpq�&�'m�}`��5[�h�c�,g��1�Ke��{�[m;���������E´ں©S:�Kve[nY���l
���*}�.���Ƌ�N$�����㙐�q�T�%���"�\�M����e*�z���� PբcT�����ኼjqX�CHT��J��dЃ��HJq���O������MM'�/��W�y*pz�����5s,�3"�sL!���)�Wt�
gT��0����A �"�������XPŊ��jg���/1M����/����_�T|�� �.
Y��-�,`L�e�(�˲)�[�0���01�m���m��n$|�A�����?�&��Eg�/�BC9�^��en�1��(��~	d��Ɨ]��� �jG�So��q��yT�}�X�d
"^��#���U>�FbjɻG!obR���֭��J*�ݜ�T�I}�lz'1���f��<P+d|!�gl2�U<@����r��x�;u����-$_�� ��LN�o�Š����iO�@��<G��^<�3�H��� ���0�r�bT��X��{��1|�+��A�;�G[5�Rj�o$�����Yo�Y1�7H6+�[/C%>|�N���hS(��]�n��;	�̤��f�������'�)}y5� G�qP�<��j��!k*@q�'���e�R1���������1Ha�F�S�A�{����^����&е��[k�C�[�QEؘ�?�(�u�A���F7�|��o���$A����n M�ZQ��ZE0��饬1^�k��M�J�#S�/���t�C�W�˗��S��� �1�5c�Z�����+`�[<��)ⵢk�%P1���E����H��$�����~_:��A�.8��ݹ��׫/ls�~�6b&�_�{���?E\O�(���7M��\�td���wPKA�s�WYn�n�^���)e`s8d�����\�8C�2�B-�̔��z��[�m�K���Q��`8��ӷ�p����`��.FsiS`�G�����`���C�8��3�u�+�	
yG�H�h���y%%�.ĉ�ֵX��	/e�-���2���|���{7	���sʣZ�G9�\'��e���p(ט�<x���#��i^���������y� �,���;&ch.��'#�4��Ew�I�I%�0��8�J1s �
�ߝ�_]_E��e�Q�[���~N�eZl��UF�N*7�	t�T�\U�����I���*�v;��;\����@c��8�2�'(�Ƀ��wU�Rp��1�&h`�sg姇�pF~����1e�e�җ� �[��4m��C�����:~k;^�l�OXM��@��f-���ު��0��_Ee�Bz�
*�9��b�D��䛧PZϤ@7psʵ�Hm��2�R�X�;(/�?�/ L��c�o&4ti���'Ĩg�k����ϭ��C?jg^�3d'�-��\��nI1������� 6.�/e̡����PG:�Z��5Cum]��]��_�*�#�.���ll�i��vL �7u�"䴠l�]���gTn𠺅��c4���B|Z��-%�H��i%�*��;�4�mG+}=�=,Ub�F~O�6h���6y^bc1��{ ʒۨhP ��`A.���̉�{���Z�sV_�?��,�87��4�*�8��]E�Ѳ�=\�nr�7S�՝`7d��LY�0r'8r�ދ�?xf@��E��jJ����N����h�yAN��"��;m���s EU��'�u&g�7z����T�R7&�n�k��kQ�tAT(q��w@ �*^&Q��.<F��!��Rﯚ.������JN�EoaEL��9�qY�K�g��������8zָ�'������t�{,�&�}�9����B^ܬ�]��@�gpG��uT��Ϸ�0�)���c8
��!na9�T �qTd�Q	��$RI?�H:q�|M��\ߦ<�)���b�U��h偶/2��^��iZ�(�	�V�B�TTX�^G���d��&�z��j^4Ʈ�0���#���I�fΠ�vY��K2����wv�1UP"�<a��'O1��Ew9je8l9��V�" R�,�T��.����,�7�L<����хw�u� XXU@t,zN�d��fzZG��F�V(<�u9[��M�2��_������8�w�4)�n���hy|�����V*� �4��q�v%ɢ"�[�J�l������������)��Kzn04&!���MT��$ K	�1�8��j���\���[}��8�Y�i�������]2�)��.���% C+��<��;�@P���=�dX��@��5�8&�R-*X�}�aF�\E`ܛBcCjϚ��]j���)Oj�L�l��xR��M���Ln��c�yvh�����~o���G(_��84�	��N�U�i�`�ާ�Ǟ�n��x�ȴ��4�L|
^%X�ȯ �Q�2O�	}}z#ص:�=Q�n�߳���Q�#�E'pR��;B\,��K�;p���bx9��ļ3(��5;���_�6#W��2�e'��)���a��jLzEI��9��m�9��d[����#l�s�ʒ7�ФAKE���f`ђ�#qBr�K��$�S��B�^g�v��qO�E��\�2@,�ٞ�����AkR���"�]1����k�Q�ɤ��Ml�J˔_I��,Xe�v��.��N���i�]x$�/��$�#ʜW���gO���o���3.����+���`�=��X����*t[(����+�=�h/��c9�#�L�&� ~������'cN~�Q�דZ�@>�m2�5�]"�PR���w+�Hئ�mݪ�P�7�BW�
�}Wi��ؽ�a�ז]���)k� e@���H}!�w���/�g��o�I�Zx���%{'���JL�ِ�K�9�u`S%|Zm�خ��������꒳��e�H���Jhe�E}��}������ wo�N��咹�����q���J+�ޯ��y`o����j�r"��5�Yg4�!TdKB�ll���M �<�]�yMF�)=�S� l�t��p2�<�:���-��g�<sL�P4A�8��v|P��&x����"�7�a��M8�|�9��4��0c_+�zV�|(��d�I�/�H�w_��c��9X�7�" ��|����K%Dd�ˑ�gT��a^�@���.������,7�ˆ�����t��j��Ul�إc�w��[�s1N�4�pa�:J$E=t�,% �]_�]5���#_���8�U�2���8 ��S�L�'!;,��-���^�7m"��mg��Y1� !�O�R}�>����\":�o.y���3�&9HX���BQcj�Ds누L{*�N^�-,���am����.�S�1�C�1*���
��'�o죜��F5�(Z��`��_fެ�-s��΂�������G?��=֋~f�/���HBV
���zq����_��s�.��#��������L
H� r�l�������6mpAm�j�f���	~�S�B�^�A�'+ռ�X
��0�<�}@d�����<��X����z�붯^C�q&ɺ\�M�B��xv�T�֓r��h�e����q�i�B�E�ѣh`F* ���!�N�S4^(� ��曂�����'����=Κ�+��+D�-cu�yY�q$M\�{"����M�E�Iփ �]�u�	�~r�!#z)@dFj-2�:$�綾~࿫�*�j��E��R�����n,�犪�O0#)�<�Q�wfy4zI�Ȃ���Ebhd�(*�K���f�
�;�8|�|;-��ەw�?�d��'۫R��+B�ŝ��n�d���"t~���mq�GkB�-_��f�$o0Sړ�x�Nn^q�!��u���8�B`�}V���r�,C#/��E_�v�g�p;)��#��ri��ઐc�p#�ِ��4z�\�j���܋����y�TY��j7$�P?S���P#�ʐ
���OA5�?���#�Mֆy�Q���S���2A���-[6�,����D�p��CU�fW��Dѧn@���ѐ��#b'+����c�"]qis�>��Z]_���X��u�fb��7��a��0��;M��Gt��hߘXq+h��)?�k�G�s�b�Pu���I2d�ͻjE�!\�:I�����W��}U�2	� W)�4��x}$�QFG��m�Ӭ�.�����U�,�~d�
+A��2�W���a%ȣ�c�8��3k�4�P��˛�0"q�cP�f�.���b�wŰ����^f`������Rџz����<�_�Xn/����i�����?.ir/�6p�	tML���˦�
�U@�	 }_u6��0}9�L6���}��H�R��+x�A��ҿ�.�5Jʈ�Ē�X�X���j6��m��
�D?�R&��T�}����1`�	�[2�2�W���s=�U�Rd�[�3�S7��(�o�ķ��|[ش�'�m������'WKb��!�Ҹt��.����[��-�>�����6���r�U�-ň��w�����u��9�Mq
)E��3&)�L�P����B[�>@b������R��&z����/n�q[k5� ,�`�b����A��>��QɺM �!/���%Y^�0f��^!�����p#t���sNG�V)����2�e-�����D���ﮮsT����8\;���\��Z���	� Y1�Bz0�}R�òF��d�+ ���e]CO4�&Ƚ�0�oZ���/��.��6: P�w���gv
1�O6D��\��ʦ��^�>����vĀ�|2����mUG�y�>%�_�|�Vճ�`��D�H��q��|Y`BYΦٛ���LZ�b%�D3�L#1����!|gj�B�k"�Dy���"�9�����bl�|b�V�.X���b�9�l����E���M��oGx;�����"�X��x�Ww�`����$5@F��U�r�7�(P ���c�W�K,W�l;_�K8m��1C��`qZ\�m��YkI��ii��%�����o{�q�A���c��5xP�Q���v��А;Eׅ�?cG�S*4�xwlUi)�C��3R��G�L���sl�V?w���@f�i��"7���6G0,����@6�x_�yM�BRѳ&�b��#�bW,�:A�?�!+´Ryx.q��35Vi�(�2��XBX��z��+��yſk�?���.�M>)(+�n����.�|��\�`��D�w>�&�Ã��q?^��%N,�	H����[A~D�m"�D�0���\�
ќ��]ڧj�5(q/�����?�.6�8��cv-���a�d?C�����U�N�C�&+��v8�ɟ���酪~��ë�[��!�8pI�
��n$�LVx���=q��V�B����S�7���&�JrMӖ��K�&���4 &�٨N��|ݙ�w_1j����҄g
�LG���`Q��<??���ho��	_<1P���?I\z7�'��.��EWۉ��|�x�(�6A��������0.[H���9�ن��1��t��8ګ^lUv�����肗�}�d�9Q\�����:�(q6R��"����a�_5�D��/�L�e ��"�IH\ K�'������x��,1p0�i9K>��m�+��m�|�����@4��Q�����_W�<�C�J4�1��nT� ��w�;�VN����u���{�O����4�*�^t�6��S���2�. ��e�R�*4�«�f���DNa�f��Z�5��@��N���E�iQ���l���<�2�၆��7�Iё�6�*,��;6�a�������6>XG�� 1>td;�����y��$�'G�jk-�5�m�L����[�����әֻ�ZˁE�!������O�?1��9��s������)��pPV�L�G!?�Gn��H���2p��f� e/�����Ck����W�	0���!Zmx������@dM8��H\fQ^����:�<[����t� �&���{d9` 9KP�O`c�|*��'��9�]q�A��[�wd�a�2 WA��KE���.���z\Ҟ*����+,��Yѐ\  BJ*��!k���H	�&O��T�,��AxE=�iǻ��"c�2P�'��N(�۷��hE�ן�p�xq��� �0��( ���!������������>p������׿��Ou;�ȅZ��Xo��H���"MSX�M�t�%w��X<���4�T�9.��6��C�li��j2ϸ�9��[%mB��$+s4�>[��'A��Ťt&9b�,����I~����yK��=,�n��1hS�x�y��_R�Sp����l�8�5��e�69x�u��_U1�-�zQ �Ԁ�^�mx��6A�!��c��e1��0��M��J�������_��ү�M��놐�W��ي8�Pwq�M��-Q;R���P�d�,5�-n�?���	�kN��d���)fc��QE�\����P�$̈�Ȝ=Լ�o��,�m�y���>�l�AAL��A�eQͯ��ޟ��"Z�C�Ô��d?. �������ɀK�&��Ly��X(��;$K�������]��j@"��X�!Y�����/0�fR�7�7&��z~̂��b�D:j���V�y@�>��<�.�X�[ՕJ�8�=�Jq}6W�M�h}�+r�mnM�Q7���7�n�DdN.n�~~$�c��s~PL�,.�ymޘ������S���&U�����|�u�����Ƣ;d��>�.�$��8��Uh��	"��7�i�[L�
,�XB����h�
��+��Ĥ���SX@�����;Du�bje�ߗ�}�����Z	ˈ��=��Xc�Ho)��KH_ȅ��o"�:��^�~� �*�(�%^�,��"R�>����Q�ch����R8�38�T��M}>�$��l��ԯ�`̤A�-���:U<����K���WrX��u�  ~3�=���`�o����';�u�p\�ͳ�m��ʘ�^T\9Oy����_�H�/�A��:U���y5f�Q�nq47U��n��׼FIBa?&r�ɾ��	��ux��h��	�r�.�?��������M� �3������D��/H\�D���,��Ti��q�Hm�`h�؈Ȟ����m��b8q�;cc-�bxhTm��Z���ži�̋Z٢6J�Yc_�Xr����:8�bI$�U��S��0�3���ž*�ת"�E�{�A�6$���"��[�D�aR~����6�[��l�ypaUr�8v.��ZX�=N�;�K�&Q��%�~;hE�����40�f##�"���U��?�0���+����	`lwI̽3������������V�7�<.J�kwm�'�d�.��Կ�����qȎ���5�1������aKo��p8��k@�dN4�QL���F%&s� �¡��?J�)��>�B+���L�۶�\M��Zu�!��$Ӯ�U�/r;�J7т�+�A�V��0���T鞜����y�T���ޘug�J�/�}͗q݇��cMW~��j-�}d����3*n�*���=9�:�M.K��H��B��8��͵�Ls.j"��r��Bw@��ڲ%}��.��!�A�xr�Р,-�o萛� ��1�B�<=2Uu� оk�!{;(�6{�?2�L:2ξ�N�㧵��}�n�3k�]���
�bjjU��U�����qw�)�g*��
6�'T�<�~�Dx�!���N��o\lS��P�fq^�����]�o$�+�����W��=���=�TqE�0���]�"g�|Q#'e��y3t�������o@��������nK��M��r�U�C\ɹ�%jhZ���� �h�Xw&tS��TOo�f�qH�Ɯ	H��&է��`׸BȬb�L`���R��b;B_f-\��x%t��|�����hHު�P�z�)b�u}���#mA�0^	?F�Ƌg����+�X�2�/�QC1y�GU�n������4�j��0��LyA�1T���R�xE�F�r$�ߔd�g�,`<���~��Zx`���!�-�T��ǆ� siS��v}"������%+��7�_Z��T�J1F�9zF6� �ۋ�}2�y�����^!Wy\�Lp���� ��۰,<xf�%�tXink����,P�Գ��^��{��c�ÏV���kB�e��g[ը��C�$�3ώ	�bW�[����vi��tvG6rm�[�$�����2�k��*��ݏs�|���q��Y��)�|��p���*�&���z�V�[xn����P!ցp�,���� 񨸒�L�^W<r��(�4�h��������49<M��>*Q�3�34�DTS Ӡd5X��^;oHٿ��gBF�0i1*�����,����-Zao��ȣI/��~u��R)���k�!�ae�q2A��.ġB��&�	ݒ�h\niB-yˉϬhE��9{��}L�ą���}+�3S���f�שa��D�e�A���hp���n�o�C�ב�����h�6�����@�}1�3R��}���	�wЊK �,TZ�}?��C��kK@�)�_�4Ҙ��  tn�k�SS"�O��{dN]H�����R�޺ �	��_�6�?[P���V$
>�,�|bX^�͛Y��T�C�4+5츛D_�0�X�䛌5*DV(`���$������E4ϟ���f�_	��W�%�,��C���e �[cϮ���6��C�f2���
�i��<���q;QY�m���B�i.�J��+F4�!�D���i�!k�#�B���w\R��0�b������$K12^.A��������%>�AF�7�i���Ⅽ����]wyr�Hc���E��a!w?)���UD
��+˽x���tO��{����y5�� �tJ>��n0,���^�M�,sTfe��e��M]���>�K���h<��8��}����b��`ZӒU7�-�ݫ�Y-���Y�Y*U�����*�pwH���޹��:e-���闗��܈{�Q�0��:J�O��=��i5-ɯ�L�o6FoC��̪���7KA(!�8�ஔ��jוT����u_��#�t���-�r�O�k��e�ަ��4ovw1����E �G��M��VR?��o��';7�e�����ʹ�a�����࣏C�q����x@`a�]�g��V�V�ԙ�)�K���͘��"ju𔣄0m�p��!�R+����e�ô�&X��1��ʼB3�V�0�K��O�:��؆��W�c�e��F��}}�\kD��qS�[�橍v��0�� B���rz����]ƀOy��ē��&M1^�F��ƫ����}���jrf���O�}��i�R�-�c �o�]-^�ޖ��~�22�͐v��7i^��5� �K�P(;G�fz���UOq�T�&��������������p��)�6�-���!2�E�d#�fv��4�K+��!yʛ���I�(ŋ.�D�+�1z����V\I����I<���l�i(A�j㍅��_'�%2׶�3�d�B~�w|H����F�妲�}zو,~�]PA����n�I�fdݬ�ږ>|�����uc]O�ª��\�����k�]N}=g9����т�>�v�|$�/Xj�Ј�;�:�M_�Q f��k��O(�=*���iS��aY���bN'��r��zݠ�2r�� �  <�zl�O�ΛƮȃg#6��!��m~�zet��I�k⡨�#;뀠gԌ���#̚(�N!��,�-�h+�7V^�;����H��h��L'v�K�9c���ɹ��
ty��á��5k��s�v��*��%�z.* �(G��us����]	
��IH�I/����	�o׋�p��U,X����C0/-��@+c��P�6�l�H�� �dEt�'Es� ����V���"c+6��?�7��5u��bL(��P���T?��ʵ(����=��V���f�n��9�&�Y���1��b�c�:Ԉ*�7+:�����I�t�H�8��A�h�7��Cn�~�k�r�Ҹ�;����d����[��й��圣'�ѝ��d+ۺI<�@�۞o`��NL���,��,]v6�-�}�+�c��益@mJoЅ���bL�Z�ʣ�;bU!m�r��Z ������-�
�j��ϭ��2�$�Z��5,\a��r�I�ur�e������\/}t�d��E��i�}u�\:ts�2@������S���_�1F0@�j������K_�[1�9��%m�|�w�����q���Ta7S}(�X����)i���_���Y�k���v�[ǽ:�#%Rx�+t�c�
�޽��%g.UzMzm��`q%��8Sb]��SX�b�*y���~HuB�Y�4=��l�k2վ�[����:�-�s"�Z�i����dG>-�ځ�iQ���8��OL�j=L�u�"�c@�^��Յ����5TI7��s�m�H��ᆼ�D�#R�Ŭ$&`���" q�9b@Z��,Zu,�bm(��l�h��CC*!PŲ�σjy��J��t�8��ϫ��r��_���Ti�8�\�y�����6�3hV�,Q�H�����
�M�ʓ��ޜף4f�%�/6�*\Eԟ�<ĉ�i���4���ג����w'"h�i>��)�������la��~L#�6����$e���خ5
����j��Q@��������<i�v��-� �&Mds�0M�J4�QU2]O!T$Z,	��ˇ��N�'	���\�9�j� CP����!{�F���}s(�6F�6�<�E�NJ��Ay��a��%!5眽!^���T��T�L*9��	bѪ��/b����qp0@�ܛ�Ќ[��t['m�{CS��5og���`��=1u�k�ʜ]��*�����x�k�b�L]�?&��s*���^��t��0!n OQ`� �D��w@�cƻ��K��Y�/JNq^N��R쪞^�|���Uv��fY|�4|��^�����W��_�kq_?���>\���f���$�+�����|������07c�����7w㩿�wl�J���əyȾR���LY�pT� b �i�'�N+ �e���E�}�J-F����ߠǍ��ޚGc`'�񯁥~Gv�.���-��A�pu�^��N��K� �L�O�j�V��-��u���@�d��"�<��(#�790׻D�G�0���oP�9�r\�fZ"}����4'�:�J啩��(�H&8�ҏ�jM���^�q��5���!f����B���ER�7���M�=6��4^�M:�/��^�D�²ง�f͑���1�<� Kj	:ä|��mW"e����w�u��	ձB��&`:Yv�=�-t��xg��w7V��T`6�Z hk6�ک�'�V���u]��M����q����}x��L���K`�÷M0���H����j����c�6�M�b��2����N��T�Y��VEt�Ƽ�&���ۥZlj`��t�l���o�]-(���R���g�I�B��C���S@%M&v�F.�FI�6���L���Eq��L-kZ���H���@f�A��IBt���Y�CU�O��p��о��}e ���.�L��J�8�9��	�a>����cױrZ��� �ְK"�gt-y��t��y��z�E�$��e�Pk�+�W�!��X_�F)T��tr�荢��tL�_M'�h�{��y	 �,��n��@�*'�I����!�pp�a}���%HD���[��)N�f���p����BN|��E�*����Ŭ��Q?��C�����M�K{���9.�C
Բ�)�F��+�i��-uO�inO'a�7%� �12�2�C"2�Q&]m���(��-z�Ae~WH�l���׊7��A��H�I0W��?0�ᵟR�S������F��?�adѝ9`��i��6Yb�䫻ĤϨ"�}!��r�4��>�Ș�����FT�:I!�a�������~<��'8(Z�Ƃ�k�JJ�~�b�?��t,R�v��6�Ӄ�?�߂hf�*�e�&s�w����yH�Җ���DU��}K���-}G�#?�/]����C�b���ƯX��G��*���T�71�q���k��qg��je]&�O4}`�˥R,�S1��E$?���O$�j��SY;Ȩ�v^��:*d���8�����8Ok�rB�Ft�����U�*�"�`|e�*��W�X��z'^߷N��kM��ǵ�"t�*;��C*]qL:o�%+.+0�� `��NH:#>����L6U�I�F�wT�IO��g�Lal6$"�8u��7n.�����[�2�n����} ��Nޤ).��Y��y��,�xi/�+�11�����b��`=���ݦR���]��ˣ�����?�	�
����� �d8�w3t|��-�_�m���u��w_�Ҹ��T���^l����o�7�.N�,��e�8V�L^d�x�#ح�&���J*;8z��w\�,��7NZ#��Z���`)�T��@MW=��wp2>ڝt�t���rŚzq���.�	@h����~]�w�_T�s��	�_�$WKG�b�4��S���A&�!;�0)չ�������N	�����WbE��s�+`e*�r��o�g�,�n��a�����>�4L�"���!�rW6�������,�Ɠ����;28s�{�3o�u�4��V����a.5�I�{�A�n�k��7�o����;X̾n&��Z����m��Sdv��ơ��v��bdu�,�@e�+gh�AK�O*�s�`����AD���&�����"���9����^�!Д6�n��A$��}�Y~�ڀX\�Q�}�u�{%�����oUoT���H���������p�|ή�}�N}�I�y3m��%�$w��"�!�IR�Fi3V�[�7�7����$����RǴ�� ��B�'�և�N��h��J�_�^ҰT�Alx�k� �*N��y��� O�&��h0"��������rP9pՊ׆��p�Sb����]�G���b�{;�����YJ���^E���I 6�xV��$�E�]��T����`�O��W��f��+�?u4h*�b�i��'7���{��������4�#\� $�-�m�\����;_��ua��[�D��d]�K��b#s'�"z��#�m�#M ����P%�l����ז5���2�f�+��%�l�3d��^l�c�A�*mR�6+A2(���P���Æ�}�d�g�����_>���!�Kw%�gv?g�������:ᾚ=�����yJ_ ?m�kL����s�8H�n�˭aۂ&-�W�*�d���VA~�4�1e��j	⫦�R���T���6o��X�rԧ"�W��i�[e�d(�=��=a��3QPH�Ϛ 0zF�R��+�fۿw����*�S���~��0�Щ��^[�r�/�@y2�(����7_��2Z�ki��$&bG!K�#~�c�����WF����^� r-،j��o�c;`�k"jM��l�f���c֡�g�/�����+��;��,*1�����+�Vm�$�f_rW���˼#uqn̷k��G�Yv�ᚁ�R��^;se�z��	4=�?�-C��c��6�C[(G��z�%���X8�9��j,���"_��j�c�E���4k���=$�>:�2�	o��(g�2|��Hܨ0�M�(��q��秃�)1҃oC4����ӫ���%���D_�O���""J�̠wW^��,ф��<o�?�� �)�2�-�6i?"f/��L�����N���S��L���x�������i�`1F��ٜ,�%ͦK�
t}+k~���\��`�e�	����H��Is+��|_����	EdЪ�� ��a�m�qك�W�C�,��g�n���CƸF�?�a�Dіx ϓ��x7�������/_��bmx-Aq�[!x�鶅�G���{���b$Քz

�
u���� ���I�6ֹj�u�l��ר�����R��|�!h�����	R6aZʦ�[���|���FA�)�����x�!S�w��w��?u�������N�4�H���c�>���<�7��ur�H_���L�p�ж����ή�E�iO�`�A���)*1X�Ѝ�����d��Z�q#�r�kS$���Ч/ørG�@۶�ڃ����i�:`+�Xc���3�~I(2�v����WT�[�Ԉ� ��VӒ!��Gi^.��ى:������A|�eF(�#�nLH�c�iS>Ј7ǔ��h��?z�Y>�]�p<����G\+Y�v�K�ߛ�w��Y@�Y�"��}D^3tc�S�M$�L�jgk���'��� ��^�_�~�؟���J!Q��l�pc&��H�+��(�w�ԑ�pf ?���n����[�X�P�A�	!0Ʃ���Zc���B�2��%������U�W>�h-�:�S�"�8/1kYyH4�xt�kg�ݡ���n+O�`��̜����/�I��\��3��<�c��;�_$�خ�={����T^.�<������>�5����W�u^��@���G�U�?X3��^y3������FS��<�i��
ˏL�j��/��i�>z��,P|=�SQ0̖Bn��<.��4J�_��O��5w��ii&��/�k|�#���z����F>��Ȟ׋F#���yH��D��6g)ZW�wq!��%�������wӈ!��c�>��a���b芰]2K T��1G;��Y�(�R���dtÖ�����?�Ȩ����X���0�����?%ؽfM��]I�s�A�b��;_B�@��^$e�_w{��~�=E쀆ߴ����m�
7��N�<�7Ӝ��S��'�%�?�� |%���h2���{G�uG:��u�(FpQ�Ђ3������	������#Gn+��{%�����C@��<��Ë�\ւfǾM����Zج�Ѽd`P�n����E=��t����Lc���������:�JN"TMGR�a���� ��V�9�!����g����2`-\�iڼ��u�g���ԣѮ���l���I:��f�~3�0e(�0���	ŀ�?)��Fr�k�ĈI�x[* ��[F#�"4��v�����^���r)��9C`���g����.�}��s���Rf~��#��\�����'��i��bn�o��̈������(ܶ�jZ(���eDCa������4Q��������mf��?';O-��1�}�#��2�K1�qת�B�x�!�S�\�)������{H4VDI㎯'�H�g��P�m)���ogR��R��g�[� �����<�B�r��p}1=#/+>����h����o�>�/�<N�4o�;e�<�XN�4`p�qٽn��}fi�i���
�W���h�Jr��W�i�m�7��槓��b�w�	s$�B
��U���v���4Z���Rk�]&w��Ǘ����*�@V�	�ǡ�8����&�{&��U���l�n��M�o	/����>V]�$'�xT&!�s��x�Y����YJɃ(m�Dޠ@Y�|��o�,
dG|N�'��L�e����g�_���G��7&�*z�af�dr�j��|0����/�_֧��m<���Eo��)���
�,�;��6�c��hTԲ�����1�ɲ���}�3"}.��f`�YAޚ�@��+l�2����аYz�H�z��!lE.���d+# ��ǩ�45��ѝG��P*4GDܑ��֘oQ�`�G����j�|��O�a[R��q�l3H���-z�6F�0�n�=��\%+�p������/.�
�0�	��hz��2軳✑<zF�$�->:#�#���l�iig���'���q���_��-\�0��y�Q����Cz~fOJ�܊�Oݜ)�\u�Q�( ᠻ��LN�&'#<�Ҟ��fKi,�~���Wp�8��1w�bQ��RU&�e�˄�Y;�h��>hco�~�P�H+M�^q^o�O @S4��-���E��v�Dg>�����Ķ�]B��4.�܃�N^Ī�]g��-�Y�����ėOS-x+��eƗ���>2��0\�A�_ ���hZ�؜��w@�]��~�z�6LÊ��Tj�����o�uog�ʧz|X�U �h8g�����>�v�j���ܕ�eL��PZa�˗��c��CjPk�%� *���+*Z��ޔw	|��6_��@���DU'U�����!y�HjXd��׺��{>,)�9�M���.zq6a�΂W�0���b��4�M�W��iR!,^�ef��n���y��0fw?�	���"{٭h7!}w] ���c��N�<#l�x.����D��nҗ�y[jF��a��X�w_X��0E�T�oX�d�Ah��rF �=�=�(=�ޥ�
pAAYK����z��uq� �S��#�q�+��1���q:��mOQn�X��b��	�eh����6� �Y��ȷ^��9�ܽ�R+�����Y�u΂=+�fc�c�tt,#$i�56��m���љ�ӎ���#i�<�'�a�>](�J}��[���^f�mѠ~p��?�d0:���;�U|`���t$ANq�sԙPJ*X��%�����c���Q���owB�IH����S�7��3��{�����~À� ��AP/�Q���'�8���wӇ�jXYc�(w�^�����Cx�,�j���~�"@'�QZ���@7i}6�O���ܲ�rR,��&�{�nbA��D���)ϜFԫQ�w"^.	��v��?��ڵ�g\l��B~&��V�w�vC��`f��Kb�p6�mc���ω��E:e���WQf�m!��l韧��pɕ����VcA�}Bh��l�I˰Q=��t����>rR �^�C�qؗ�qT���:�r�*�F���L�Vl՛��Nх�� �g�Z4�aL�g/@��l!�H����;T��g�zi7�Zw��U�A�4�L\�C�#3/�R�
���"�L�ʯ��QH�`n]7�y�U�qyb��u��㾀��u��M/o�K��R�q�h+,�F먳{rBь�RZ�s�]�����V�$G��1�*���n%���P�kl���!�W�C�n�B^�/�׹Ǜrh@�H7R2�v��E���M(-�x��?��L�H{�g^b'����ܪ^q�
~Пɸ��	�5�����.����q� x��G��{ҝWIN1]h��-�d�=�R$����n/�&VB0�n1�Nˀ��2�N����y}d'��d�Ov������S|cz?%��44/�� f9��NqR>�n�נ}�'�),��f]�y�����k�bU%G�h�9��gwj������J�nXI��� �e��n��Eh���R���س�mL������<dsA�����@�Ҩ���>���`���-/S�����x��	��#�Q�\�Q���Vu?�/!���P͒��.���?P��Ws,v����]�͛�h���H��%>��<,C�C^M���~}2�
�h3��,`	/rxJ��o�ȧ�vE�D�
�}/�b���>`pC̝Q��tB/�k�����`����y��:��9u�H��'ޙ�!�&)�ؘ����� A�����\Z_A<��F:���u�n�Va��C������8�B��A%�b�-U�)��R��L�'c����Í%�)�f��ټ|x�8q��f�W,�5 ����K��!Ed��x��1�ht�ٽ�::��L����º}C/T;>����+]�$nI�md�܁���Lh��1~��:�*e�ʩ!3�o*�����������h�&�E9
)����q�%&�j�{�x��1�ƹ�<q���v�*����f��M�!�1�MEi�d��9'�����%�n�7��(����'eG\�,�4��"�n�5Ź�ZJ	���<�Er�V�R���k��.w��gf����<���i�@�[K��T��b [��t����ܾ��ܴ{�f�*&Y�ʀE�A�!ʬ�E�����Iv����x���%�%�Hb�'�������O�_��9K��09K�}��6jJ\�����{+T� ��wsڤ��c_�P%��.ӵ�?E��ᾖ)a�hmܒ��HL��1#�T��X�4�/4/��V����> UI� ����+v׾ʞ͠��8�}�!�E޲l(�����]x)�Ǎ7齝 m"<�Ɠ\-/5O^u�A����E�0S,GB��2S���h�;_�=B0�>I����[H��
Օ�R�,�����m|��\��Ύ`6%�k_NT�$/��[$7Y���M�[�+�0����4I~3�V2����)�/Ls�M�R���y�}�[.�[W��?>��	��������>!�x���Ӄ�ѝ���l��r����� ���G	�i��^�~��^U���{c���ʊli�.�U'9���@���|�1�U5�������f�6 iO|�6u<�I>�HG���-��2Ōʳ�ng�	)��p,O�gv�~b��:�I1���z�Rq�Ϣ!qk�7M�wV���]/�B�"zڍ�.����EX�N^�W�S����f�8oJ��t�[�OD�?e���آ�v�	.y��U�0�ߧ���K�=�e��	sҮ����xz����tk{��!O�ʰ:��d�$�D;1��ͬ��dF-�qA�����*@ �v;��:��Ӌ�%FP��8����){��L
��Ѣ"QF��&��� ��*�[���q_��El����Q���+�i�K�
h�n�s�s��dE|ba��gcm��32p��Bz�� x��i��S����s�����n9ȗ�HH�ۄބC�$%�3��WSN���b��b��:opN8F��Q��W}U]*c�j׿˾4�O�Wa";J��:�6��rH!���x�8ei}�\É[�-���	Rz"�I�Q�\v>��-�[���i��M�y,w��� {$�fvA�ǬuU	*�o���D�'.jZ�|��G[�V��3e�j:�=]���щM��t<��/��b��NYЛB��k���Tɉ��֩?�l��Ў�gqw$���2�qV]Z��Vz�<��=�� ����~�g����N�?���~� T���b�W%S �α��-�X��,2*�����g��Z���McY|�D�bt���.ӽ������l���i^]\>	'A,b>k��pO|
ޭ6�y�64������z&3cg�'x:"p�U��mݘ��+���o.H�;\�����We��>�T�X�����Ly�/�1��4%O�,������C����IJ�{��h^�MD]�X��&C��bX�6��tְdL��D��������O�d�����BE7�(1i�:v�3�/zik�mu�U>������}|H���}�$yv�BA�R���O�kOW�/���&D|�`g�BvYO����!�X�Q�ד��S�+k88\�V����T�FI�%�	���g�
d�bG�'��=�u��s�]l��|7�D�X�w쒍9렣���Z��?�M��ay�[bJ�"$�� gF���_�XjMji���)�nW��&#(����l�&;��=��h�wǔ�煓�0�p@@*�d
��S�.�2�T&�0f�}##S��k��p�9�����C�HH��qr��?��U�B��f"�ށtAHlfZR�+�H��)C�?��z��<wK7H�OY﫩8H\m�RV\�)��B9�iM�{�/�eҝ�3�_����òM�3cO���*�����i6_�t	�t����y�h_��x���k
UG���}
�,۾fk��`��k��@m4N�Keެ9p����q\a�B���a*�G���n4��p�?�`�3��� crC���
�[�A:��ϭ�!>�m�@��y��R�Z�d5^Tpn^�n�2�`{�'HX�҄MP�!�S9DĈ��j���0~�����ד���.�D�Bv%�=zKXme&��܋?jo#�C�C�)N����F� v�~s��d{���T�٪��;��w����W��@%�E撸u�I;;����"H�W=b�ʣ�^�Ѝ�J����ω�/@'m��;\��L�H1~����͛�$�'h��=�C4�i�y	��h�?�>�N	����i��\�t�Ve�I�g�I����-�3�in�%(x�76�Z���:kO��
/�i0n�h�Xc��>�(8b�o���E�N���������،WxԢ.�j���~�|S�s���=��s��Ŵ�Q�9س����ǈg
�2�}8[������)�[����ɾM���o��l@M
|��ד+�礙��I�@��}�0]·�S���ƑN@,�76�`V ��rfؘ�����x2�S�`%S�a���o{R��,ݤ�c�:�q�/�Ti�dc��~�����ӏã_NzT7��A�s����M����q�	!�ݝ���utܿ�Ϯy~M�����ں�ʕ}��w�����>]���j��CT��nc�E�p�1��0�&o����[�n�W�n$W���t��t���_����˅�'�
�� Y=o�w�&#XOe���7�\�hL�f�=���=���bG�4��}� --z�z`���x�&���J=G�`p��z�= �T��(;;2I������)z����C��&{^&v�մ7�x�dI��)��cm2��J���v�4U�����x3{���Y�R\���8D�[ԑ?��~�ZQܹ{O��;�P�q��|$�%�]�Our���g������n���桥�'�~�������D	E�jU�O5R�m��b҇�B�
��l?��k�φ���/Ñ�vJ�ܹx�;h��;~�*�}/��P��|�Βu�Ů�/0��{�W�fۈb��2O,Yw�&�(R%�� >��;�ps��K�r�`0�;L+�I��J�|��1]@}���( ��-hG�頳��W^	L��X�U�A�:�K:�I�����AE��C���(���h�W�Yzˌ˅�z���F�Io
���c	`! ��e`T&�}A�ИHOç�K�ŕ�����f�u������_0�3*�v���1���I�xո���~$�P����p�;��>n�X�N�1I�C��E,���z���.�ϭ

���O��[m�[1�Eu�$T�-���h�-��d,�3�������k@��f?�ޜtP�Ygy\��K���g)l�t�d ��4z4�I���������x��F�[��c�[N�����~}�|���"��=r�
�W~xȍ�����E-&�q�{bA�t�q�⠶�mu��q�1
�s�;+�צ##:<x���.@B��G�c�����{��^;;�N�&3����8��~���"�սЊ������IN�|�g���-'���*��M}�����<�
t�Q�Y�+U��L�L�$LV��y}!����y�#�k�G�\O�^g����<_�cBjl��=w��^`-G;�UX/I�B�z\^~{�`��c����T��<����[�\P�1u����TM�6H��)���m�K�����͠��'b��8C��g�Scƴ94#��WZ$A\i�jΎ��P*`���5������w*�v�Of���n%�/-_}��L�X{?�_9ncH��,(��gO���7�#�ї���	���~���<Hj��������b���� ��^R�THE�����!'� Z�Bv��Ӗ�b�YL�ν��C�ܘ���q {�e��f&��p�IF�����
w����]����ui��<�+�4���8�+[؏�w��9��f�!w�à���@<�1x����B�%���-C���AZ����N�M�����)M:�Q+��t	�)��烿pY+K�%��Z���b���6P��Q�)�����L|_A�e���S|������,��s%b��W���N7d�,�z�<�,��Ǹ��h&U7b�x���&�hS�����}�*�������C��ip����u��#���'mU��(p�����z�]�F�0�O75� �,���A$����S�.��&{��FLF9$ܥ���;gH�n|��sZ r�sqh|�Z˭}�0ѻS�[E�ljM
��Ah�M�c�c����.�����S[ 8<AM�4+ ��m{Q��*Gj��N,���!�5�u�J�����-v�P����z1�JY� ؞�l���~.v��S) �둌oe�l���a 9G������M)5�綥ll=D6l)�AF�!����������#����&,30�,�Kt������7�vT��t���srB�zxz�<
�3]2��;�]�����(�#���ܱ߻���srI��D�5�>�6�����F��ӓzW�G~z��-���Sa�������)m�H��K~0���N��M����O��T٥�FTn�g���9)-*����iIn��9ˆ����w�.�pՎ��&R5%����Թ��P�)�4�W��^J�!�V�L�Uz��ްv }�1��``�80��S^q����U$�����|��~]qT=8:�p�P(� x9��������G��}�$�YG/s��A��4�>Lہ�u2�6�H�����,~�/�k4�q`{�r�;�'���?����D��6;����]݉y�']^��N�$AY��N^?�@�=V�@c�J�S���:J�p��5)��M�����-���ؾT'(D�O�-W�Y����Xϐ�\�A{6 �u!����h�D\�����MX�ݽ��t��aq\ R��d�u�-���TsK���gD�����ѷ:�Q����g���E��pߣpH�^v3Rj,S}�b �.X
���N��Wܴy�Ÿ�bL_ǽ�Q�H{�p��/�R� ��~���5؎�k�}�C��-��!�ȇo=kK�5�%� *�0}����I�3}�8�S�<���5ʡ�Μs �1m�m�R%��)*�*E�l6�ܮ�q;�� ��عu$����#��^���-/����A��;t�NB�}so�+�]��v^�v ����i��/!Z>�K����-{�C��f� �M��>d��y�RJ�S1%���k�ۢP�
n��U���E_7�5�G�:��&�� #E�]P"I�����©��������[�J].�@�-+t�V�F�*rܩ��ys�z�;�^�29.�,�F�{��%<�a��'\�����,�����������jJ��EI_O0���{ȡ���d������"�������y�4u��
�o�� ���,�#[�΅���'�Ff����³�Qi`�����6�SD��n.z���$8r���`��XF!iؿ0a��N��2�^�ٚ���.��j��,7�ل)>k��`eҟjNt�����K8(��'�	�١�V�g��IC5$�Xp��԰A˝�+���K�#�s�o�*|�.68�i�����J���F	@�3�J��p�`��IE�4\:�F~���5���8���!��J�et�;,��$��%!���̄�[[�)�?��kob��U����d�-w��ex�W���k�WBٜ�m�2%�\{QEϺ��,��t���C��}�|*?����1�A��pTϳS�@vPB��\�2Y*�Z���1���ڙC��yaz"h�p�G��]�}��1�4X�_$�.H-�Ռ���d>�鈫:�V��֫v׬��Ae_�wYCwxou攑dwj�Pp�VM���ۍZ�"U�,�@5�c��w��n*̗C�7=-,M!`=��ζP��ʽ>�N#���_p�x�<�z���G?��^��j�-�f�3�K;Su3KzA��΢���Z��z��4�cwC_�IM����R��g�^Au��	X�wӈ��wֽ�miJ)��	�ESSL*�rh(��9$/je�q�"�Xr��i����9ۧ�RN���,y��}���n��i�� :(�5�j�;{�+�x/�Ԫ�&�ڼQHP��/����Z.�yf掍��5Z#���W��x����G����������Ù�T=v\L���$o�/��v<,��ȯ2D�'<2X�V��`]ؠ���}9m_:3z�x��� ���
M d8�d�[l��5-���cۖ�T0kљ�b8�����By�9���v�y�i�^�Vɶ}�n��[,
+r`_l�#�}���#Lƚi�C����ǯ�jG�/O�<A��ʳQJ�'֮Cz�AL��$ˮ���u�|N�X�(aV���f��P�J4��3
�$]�N�]x��|�Z��S�\�<�hl�0>�AIA?�
jT���N{t �������=9��wO3����*[�b������)M��Z�\�#���:��3ܠ�J��]k޸�I6�E:;��ULGȐz`A�˓봖	�|׌�7�۰��U�[D�Vo{	���5�E?�n ��$*���,�v	�j����	���y�P
d~LBۥ���f)�έ@���U�U�0���6zW*�����]toh���!�B�z�a�W�����Jrn���J�P�׬�5��ж<[K�@�;r�䳤*�F��v|���2�K�Pgȫ�qfldnPsSea������]d��04�N���g�]NG�J�3��U�`8b��ppm�h
�'���ǃ������bq@�e�������ZN��he=։ n+ϕ�]�Q�h�ml��kţ���#?�輲?��]� Z�ɩh��dF�bl䀥/7Q�t�l��<���d��IS&k�A�w���x��Ҧ�L��g�$x�#Eɒ��Y*��愮[���=�	5����aq�*�����3@�����Oӏ�<� ���9��s�2�O������2+�:4EJ�Sp�pI ���=�k�מ�m�ߢ4�Ɩ�+t$�0A�zР�sa�@�c4~�Ӵw�h���l�E>�?��G�2�t��\j6�_6>�9��X� B�y��K= ����(M/��Z�E�QYg<_,�������J����A��9e�Y����(����.>���H`/b�Z�����Q �=��g�#)�#=(�Z���C�F��\n0z�S��%{\���=�ɩ}.��\��O�`�j��ո��@�,��փ��q��Z�i��A�c��{ �-�yt���#���B�&��"E�Ö���|�j�W�2�g��ʄ#������G�ҊY�C{
��аr����������6�ugr��m��B��~����E s�`����'h~���	�
�>����k�ň��B����F����;�>Q�~�+O���&�e8������o�DH�����1_�|���G�	-T�}A�v�f�Mi���A3�S���e�E�0VL�N���*�8*�5=�Bknp��~�w��Y��cо]�"�ĝ)b�N|?h����h��i���d�:P.<�|g�1���*L�݁��zn��k&n�֫�pz�S�p6�JI�B9�?� �/A��j2�u�-[������HF{^�Kv�aD�Cm��笂V��YJz;Jl�.bb�S�v��2R=��[�So8�h1o��Ҡw֦���C���8��ꠜ@��xB�x�I�I�
���[.�H瑀��A�_!�]ev	�0��m��dz�׻�(��';���U�[��(L�g����R�s�h�3&��VX�L�5YWB�&<Y�I9��f>2go�Pj�Z9 +�9`1$�'c�-A�y���$�I�PZ�x��B�$f������@Ա�
��Z���1O/��.�%4x?�="�v������Sf�pG]���P��A��.zbkQ,��D.2_��t$�Y�/�zR^��kp��؁�݉\�W]�U<�� 8�~e,����|4`�]�"�-�!�u|q���8c��/��$�#��7�<��i�|�⩱�vX��A��q��t3��FÞ�҈�*�]�q��r�P7*٩�n#�l�6��1'֡��������b�n ~�C-�h���}
��=�vh�oXx嶖�]f�|�Sb����NX�&��ƈ�j���`sp�9� �6��r�K�-�.rC�t��}��gƋ�tI�]Z�l!7�S�`(&�h�v�ʳI�Z� �^���7(,3k˱��,���k��)�m$���Ja����H�E�x	9S��}��H�ӊ5Mn��0�ǩ;G�H�ՎfiM�,��e$��c�̥�����ͪ<f�΃��ajvk�a�I��yZ���eOn����tG�p90d'.$�J�4��Sxe��}-�3w�8�*�'�v������7�V�)z�l�6��Hx�D��M�b?���y3�}�<������b���Dx��|��91Z���ݎ>GWe�-�0FbleK Sgs��f>������ ��a��qݖΥ�]5#��\W�g~Wi�&�}�a��B{Ͻ#��j�5�6ɛ#a�Nu �<������2�6�l��bx1_��j�p��y�S�y]����1�d�/+���&b��@��7��^���K��n������E�l�Di��~�8w����%H��J�~5aWK��` �ٯPl�E��g��(�)/�2�g��o��?�m�ǙS��eT�����,J[_ �oˇ Qv����5@gT�Y��Ӭ� �$iD��N-Q��&?s��@�Ш��U<fza�U��Q�-����塭�rJۊ2JD���٬d���<�� RS�s��(zPs�)���#��\�{&"��
\9Hu���<�Wc���x�,igZ'XA����ʳ�L@��q6l�h�>���ſd@1
9�0����]�^+3 
�s�䘦�	�.UҞ���$m�_����� :��y��T#�E�|@@������Bj͚J�DNg�ƃ�,T�YU���gʚB��??�N�׏��$A�z�uh���Xⴴp4J{s4$1H�P��D!@Y/�~���:욳%7��dD})}�WU��c4g>Sz*��ի$�ф�9�GX��<]���B9�'����N���ۙ]�Pz<�]��$f�b�g�AD�p�I�l�S�2lk�)��;fﵫ�i����N�N^Vԍ=��*ߌ};oA��u+�=�n��Y
�﵀��=_;�mC�A(�I��s���S���ejM��]���|҆��I��H:	���4�w=�etS�,�S�����ml#�3�jۮ�m�<,�-�)�Ũ[��9P�AhB�g↩�R��FF�~݁T�;�V=$d�D���b��\P'����nɸyvg?��dSLx����+�ݏ��#<�d*�#�i�w23�����t�T��"���T-3��E@�D�����hl9%i*y��:M+����=���U)����J��e+p�ǰ���?���n6�@��`8�I�tg���1ג]=F/HmZݍ�)-YA
{㩔� V�O���C�#^C=�.������=qv��(#��h�3Ѩ%�����#D�L�@�BO7��4@���6��E��Yf��J���S+8��ι���Je�_�]�Û_5]N�쾵��t9�k�N!�z�����0e�k9��� '�~�� �
��V���ŧBh��]L��	z[�P�y�dǚK��Nh����,�5���}j�w���ᒀEET<4��ڭ�&"9����P"=�FC��I%�jaِ�����Bw=Րb���ֶ:6"�gi�g7��k�_�{�Aә���L�A�g���s!����`©�}�է�&�'al���s��Ղ�[ۚw��L��q���[��� ��d����'qٌ��7o����2���F�5��Da���6�>C#p�i��{���\�1���/�3,�Y�s�+��7���K�	� 7���a�Y��^k|��x��2�����i'�-�'$E�>�ϦJ����-vE��0���^K?�WX�rDc�s��ݥ�JQ}�S�/P�!�Լ�3��$,dҏ��=S���'�T��r�)����d5$d������E�6�g���+�[�Q=j�+�u�ieg� E9c�
���}
�_b��!��[��˅Y?f2BQ�3��̳K'8��b�y�����#J��GyD�E�T�m}��<��ÿ���#�20;�թ���?3��a�H�x��^��H2��yH�_G���K��˝����(̝���C �i��lݻ�n��Gq�/Zx��GK�}��$���WʒB�|r}�����Y����(KI������ܤ�!�y�ij�3b�
���L:`v\�ƥ�HHN��8��"���B����D���?{f\�QѼ�\�(L�F[�;iFm+{!@`7 gt���.4�a��[������uh��k���@�Ĥc:�{�,�X���[��g��?����v��\5��:F�FxgE�lil��)�[
rҥ�僊��G'���9�p����J����RŐR�-������A�~�>��'2����I�@���̳�SLԻ%i$!��o��i �^�6�����9��KC��S�%�p`�M�sɝb�e��7k�v�������q�$\�Q�S��V9A�{���\�����ER4\����	����ͬ���k��L͉}9�ft������t���n�+�@X��'-kB���H���Υy���'����q��$�"���~D���l�ѯ������蚒5���:�7����tNB�f]��&������@����5eJy@:�BK�
�|k_��˴��7T��!4��$SH�yw(G1-��*qC�����Ծ��hP�d92���{GL��ڟ��y@(�i����P_�G��-�~�TvՎ7h�8$�d&2�
�bַ ��$h�]م��0B����9�֝��jr�|�*Oq��ӧo`9F�}A�ا[��2�L[vj��䰭PE����� F��9;���R�6T��Gcѹ,��0�Y��5��%;�U��'Z�{���KY�S�M욊1�b[�H]3`F��	��5�2d� 3�>����:K��O��.$��B�b���n��
u�I�}����_M��;��X���b(uCu!���h2Sذ8s%qg�ǣb�lN���qS������A%���L���"}p�g�dE$��#|����]I�oد@�ȗ���K.d���b7���K,�D�W ~9Q����,@Fd>��!ĖK�/Z��3�����@�!�v��C�w	~>�]g���ګ��$A�7��!���1�b�G��Pv�݀�*�:7f@J��'eP8]賻��b\�M����6s�}Z̒��Pv�����寤���3�t-&�\#���	I� �:Mf������T]��IS7�/��H�HV��ݟ�q43��iS}Ufs ,4N��y�}�>��gZm|-�.�7�<u�C����)�ҷ8W�P2FvS/��FTW�`�������[u�R��<%&[�].[طr�h�ѵr.�A�����H�����@
��	�T�|��N�����кODj���']S����r>�$n"�:�
?�"|��F(��Аe�Bm��J�d@��P{���mo�Ӭ�Ǐ��%;�=���1ɧv��^kQ��n�|�`@�4�`4%��� $D��nޖ�Y��bS�[ ;h(G��.V�~�yt=x�8�ڷ�*�y����4c
9��z���������5�E��@�l�O��sM�>��'me�8���z/Y2�,��8�1gB�[Ѓ=��5h�]E|k1D��CG��U�%��8����NAwa�·j�	}�$ϛ��*���@c_3]�10YB<>���K��g�Sᓧ�i�|M��1?^��u����L)�p��k~ĝ��90�� ��q�t�\���|���c�D�{�IB^��M\�݂�r�=��֩��pN�V�j4y�3����?���5�b��9}3����V�?�`s�4���_v-��)fğ�ۘgr._�;���$ ���fp&�%h}���>@��NC��E�cJ�v%]��h6\Ck"q��IO!/	�Դ(���2���Z#����Vrr% )�-&	p������%c�5J}�-�k���dqn��ĳ�l[z������3��I�mm�P��FO��	����D�0�ұ�
|#��>����0W�Ve��Ō_@�urp.�4�]|a��M�������~��B���wZ��z>��{S߹B-C���)+d�U�vTWI0��!3��Y�eRf*B�>�3��J����0���L���p��|���ˈCb�
0��"j^�܊¢e�C�������6W5a	�Pr��.R���ȏm��@�0g�@	��2-�DfK�=5�[�l<�	f�8��X���S^�>�L_,���\пk
f wB�y(��/$�=	�h�)z���^/�l�AU��P$1vƾ=�������N�']Mؤ�΁6��I!������vL!H޳��y��{�ā.��޾�˞���:n0��i�Aa��}��Z�"^Z���c=?@�@�T�F�CH-yo���9x�s'A{T��/ �:J(qD�J��-)��7�R�;���{��ϖ}�i�҄�4J0cp�j\@����*�J�cԥH�m#�c��]�I"��(��w�y�#��s�6��@�@�d�"֪=!_l�0�a��[8V�^l���ǧ#�uf��F�?!w�7���*{Ԕ�1sn�9De�q�ѝ�f���پ&�3r狝b��eZ���٘�o(��|1!�΀%�"�ͻ>58��3��J���MO���Ɔ��á�%��Sq�fՎM�N���و�!n�֑`�)�֓��z��h_V���n#JGS �J�V;��ƈ����>�/��t�K�ʛ�bWj�ஶ��]���qØ�q����6k5{�@v
'���e$2s�_�xoH���N�e��y}�6F\|���%����N�,˫�u�Ȫ�q��pD�"2l&1*��*�O��tKV�9o�A���c�x��x�NW��)q����ն��=��M�d:���ڌM�"��e��������)x����o�d�T_�P�D�Op*""��T	��?/�m�,��R#9�\��6Bb{[b8� ���x��;��z���A�5����
�)6�m�=���$�tUv6�����>8��w����y�8���S���E�A϶ޙ�f��EC̼/���ƧG,���f�y�m���o\0�/" ������Ϗ�^�X����&���D06�m(c���F��m;��S4T����:�6_ �1�֏�`�4<�n|��Ԯ���(^�f|�Y�BS�Nd���W�rKܪ�+{t�r�
�����ֳC�����K	���z�+���E����[�Iv��?_�M� ��?��O�g"�sM|nj���R�H�oH�q7ž �#ɦ��BF�{�߰�{����ZaH�&&m����jQ�J��t|?>�w�= {�e�O�'ZiW�?e�-!|��S��3@�/����A�rbD���l��l�F#��#|��H$�<�tc�$D|Ry�\BG��A
�ڄ8���1����!A��B5��Ol����	5ttUM���@�p�-W��t��AC` c��9�4���z�G�aǺgR?ʫ�?�r��2��/
:K���S��)C�^|�F@�l°����V�n�o��R6���ѕ[���H���(4�*slI�[Y�>"��WQ�q
k�S�O���q#��3P�2���4��#u�GZlɑ��2C�@Ǆc��x$�v{F�2�q.�ߠ˶�O�������$`W�H��-�[L�_5j�G����b�G�2����w���=[�T_EM�Y��æ*L��|2��R�	%�zy�r����B���ڹ1��୮9���D��R&o68+�ȳ�-��N�9�I�|�lnqb�013L�z�����N��������A�-F�JV6�܄CV��c�O�R�&�d�lK�_o�X �@�(и���?|5�j�.�I�V��D����=���_
-�����}���̜���C0Ѓ ~�
���Rѳa��*��w���oׂ2�-�LM^L��e}�R>a�^���C~/���*	:���7���J�C0�Χ���r�Vר��`���Ja������{ClSr�w$�{ٙ
;_��`h��Ya{��ΐ7nNW�}`�*1I7&.�[�5�>G~����i�قv��O����~Q�����Z�zi	C�6:�cЅF�~���%6g8�� �*��vTe�^	GU�-i��AN�>�g*���S��k����U5���:0�vÎ!F���&��3O���� �ʔu��j�H�����I/��9кKr"8>"xb�������20�)��?�<��tZ�0AD�����M@��V`��Fvq� ��nB�4���)~���kĪ�.rx_˽�N�IǢ���U�C��6~�V�w�}a��>:����U}����M�.o���c�_�Z����j�~�P�@E�H�D�QD�$�2YDBQ�_�7�����*���UV�{D��v���Z����Ƭ��x�J��\"D=�n5��(w�ꁻ����@H1�jhY�+�*���"YC��$I	
A%A{���#��$�-r�B�#=�5}�+4�A`.+|;p���b��$6���N���)�����>�+ɽ�����A�y��T��W�쭓�z�-?���~F@�H4#|M-MR/3l�S�K
�g��M�S����"*5�V��L��F���3ȑ㟀{?�h�!�d�Ry~ ���x�IC��L��1�^%���S��j�
sj�qDOm�n�&@��9��}Po�%2!�3������T�D�/���jJrd�w5�ez�u)�qa/G ��FQ�+4E��!m����rь���Ԏr�~�ȱ(�#}����,��Jk���E�T�­�$C��d�O��8�a��ރ>�V��<�䓩f_�F�\��[8�����}_��DϬ��X:�cݟ� �3�G�6�ءV�4�R�\$� �������<hA��u������o:C����T(�҃a&ם.��~qm�|�LE�R`��YC��������d�
��K�Q\��x�f�''���Oo6���.B@�AXɪ�$p�*jxL�$%ՌU��ie�s8fπ3qf��J���-�� ������~}7Ol\2��x�dg�0T�,�玸eDܒ��*Ku�~����ӬG�j�%ޣE��B��U��B:���r3q��hb�׌�ؔ����Ձ���Y�{лuiT�zPX,�hF2�ئ�v�b�&��HX�;� 
S�y�K+]q"Y]?� Xc0q��r��� �l�k�CU�7��M�jfy*�)����I-����NIj������5�/�`���c2�4!�sAR}�`��.l�w�
ބ�"z�,���I�����5g�+'"t�ubOH��+�����gI�>@�U$<N��CU.���V�M�*8ZAi��:�׾)x�@��n~�v�{���2S*0�}
�h�b# [��/xW����gc;���z�(޹��|�?3����[b>�f"qƍ����>?��6�Aɻ��y�`,֢7��'a�J����TT�����͏�_���_��iR��B�KO2�,�����\�V[�k
�䜔�c��ep��TK��|G�����d9}s>y�o.�A���i1�����R�l�4�P셤A��������S��ga�z�s+ͧ"��g�X��jՈZ,��v
��������L:*��i�	��	���LZ y;""�e�2���-Ti�'lP�7��1T�}W7_�Ex({�Q+݇���Tp�w�[8	Z���Y�?k���ѳh�"��ޠN�s�:6���Lf��=M���%�C���Cn�c{�����N�9��.�F?�Լ�<��+�	q@�S:��}hr��|BmT�h��+�J2#sw[��� /�-I�6>� ]ҳ-t͖Z�IR`mo['�a	G�`�cn]�:4+�&6��Jc@�\���ծ7Z>ʁ� E�&�����g���Vz���� vG�f'��  ����v?�p��������\9�o����s^ ������Y�u�xO�����G������a*ƶ�Ԛ<�G�x�7xD��E>�C���"m����J.����˃&��*�yk��X��6���K�%��PT���O���p��fz�tʚ6��!ݶ�!���)y����#���Hf�g*���2f-�|�D�; ��;,b�ͨ�P����X76~:r�N<�sbt���@J:�U�K_v��2X�v��[I��,[+�ƾ��^.��muXc���#I����4D�J�)����4䋕����`�{�����Ja��X�5�	�.}�GR��R[������oeR��iK���m���%�fO��K�i42so���|K��y����{odDl��G�r��K�D.מpǶ���>����~����Wp�uX�-�M��0.�e8�4X��ܸN>�h�~M�E�Fuj:�I+��6y�l�[�ǅzR�"��y�r�'�ż�ֳOE�V_, %Qr�])�f�GҔa�h�O�x�?@�[�wb�n�'�Z;����Z6�(��6NY=����A*Tv���Rp2��a���zGY��NK9��EƠU �+b���E��t�7ơ� gY����K��4�����֟��n�N�B8��|�A��cܐ{���5�H�o�[��x��GE�������6�}&94����td�V�	V9�E�YȜ6q�?R�W�.�����"���t׮�G}x���ʀ���≿A�������$��]����wo�8�^� bޜ�
8W�r!�Q��vD��#w�����[��-�~<Q�����w�B��b�ߛ� Wb�~��!�3<6�;���v ��%7aH�3l7��^��az��XBS��<$���H�z�p8�5s�P3���
��K+���w$WF#a�Q��H��&�(=�5p�&i�K���eG�Tr���,��z U�4�3M;��p��˲o1����W�I���L��S�1��'mȨ�L|��fV�7�7`'X�F{pp�A���5u�z��4r\�eR��̠uS0/��;��vG�e��yWv��i|%~���0]���]R�.I\R������s@V�@��L_�U^9���Ŋ>\,���r���Bł���1�3�]�be5% ���hTw2Zd6Y"$ulJJg8mt��"��K�Ia�|ܧ[�;H�v2�2�$����*��+"/��ևǽ�i�9N񏠝w�����	��&�Q��<�<�X��-~�ep�S�8��
���[�x�Zjױ{NKM���,��υ���R�?"p�F��6-��X�U���,�(����4yb�T
E��F���4d	�2ү��Q���p7Q�a�ju��Y
m5�J���$Q���Gm�
�k����,?x�Kj�|�9��V� &�E��,r��8.�ߜwzP6g�fM�X�rA�^�^pГ��)������4�p�~��E!��_����Z�
�U���}t���=����W���"�>�uFfüX�a���gJ�����
L������;�'���}�p*��`]o���������} {�����K��;��T?����z�����r�l�S��S!�!���W� ��F��n�y�ӁZv�[�����t�����Z2t"^��@'q(5�rl7�w*X��9�^O������?A��ZuїV�>g&��4*�r��'w�­-R�2���4��w��,ɾ�%s�9�x�!�$�S��F�M�&}����͉נ7�#o7$G�j���Z���e�C̃C�D4s�ܙ��`#��٬|���,��v�y�#V"�<*:'�k[�F��d�5���z5�9iq�A����Pb�]�ñ*�Z� O�v�=�d܈�,�Qc�f.o�f�ͤ�%�B�YbOH��A�����$�;-��wG�n|9j�Mp�3���L]�K떔S�wv�qL����,<W��M�g�� ��I���M!�~|�u���q�ć7�{���k�#2�� �xX2�	�E
 @�*,u� ����(�McQ�d(N�t�<L������Ff�$&?U\`��fa�;j�<��(����&��*�x���c�x������~�5��O�iڏJwk���I�9M��c�+����l6�4|f�Xq��*�*�:�M~��j�Ф�~�i U��H䛸h�F�����E+~-�2㉖�0�#~��%��,3�����`�^�3���w������P��K�_|���V9aHT-)���y�f�@��vl3�Xer#�j������t�ȿd��_f���{���s>���4/I�2*pݱ�_f6�$H7�r�amq�6�)����;;R�<)��ʡB�j5�p�
�CS��d3�Bc~���v��R�o����J���:p<$��z5"H#lZ�_J�܆Ӯ�m=z��,�Uߚt,	`�\ I.�^w�{�Y�U�\�uyֵd��^��=5�h(�D�B�[3���X`��l7v�{��Ul���"�q�֡;�aa�"�.U�C�n&0�b��.r]DM��S��ɧ�a�UxcZ@���yZY�s��
�!����1z�_� ����w�v�V^w%ҩ�A&{���Ka):h�a4��=v�xhg�:�R���[X��Ӏ�*�B�j�J����
^����}/�pC��@���1an(YVI�լ��H��z�R�B�i��	�ӄ*�6} G�p�Q]g�QY�π�6��Xg��\Z�.������A��ǲ�\Q	:����}��`�3b��(F��|�U�V�G)Dr��$]m+�T��j�,�_���RHr$b�U���"5����,ڡ!�ȅ�KPg�M�d�Bdn�0]��"���1P)����Hgۻ~/��m?��t�]��Mܳ��ǋ���:�]
C�y(x���������@�1��!�ߌ0��4��m�a�<����RL�Dq:��hb�Y���̓�̮e[�"�(��v��ҿ�?3~n�����5b�����s+�I4�3��_k#o\�$؛�V(H#���v؛I`�LS��������rޙ#�N�.�T�`�Q��a��D�dђ�R��%�h@EPn��~��>�کi�$�q=(z���&�,Y|��p9�!�`��%��[T��b8�u�aC��c�gHk[{�p��@�[�|�S������o���^T=�	B��4 �K�<J`������W+l�eʰ��h:"Ѷ����y)A��E�ӅD|���{Aa��j�s�FWH8���.�a��EJ��ECXُ�]U�ۉdA}�"���yb�r�#�¿r�@�9�8���#㶉�8k�Q���������=O> �ץwyC�V��֤�K4	u��(�}��ak����!b�o�]���
 ?#)���i�i1WW���843R(pk\%���)�BgUl �}Ɨ�>�?����L+^��q��?���Q��^NI	��2��G;��H=�e����)���t: w}�+$*Sw['�"�+��v�!j��������N'�h\l��ђ�Y�r��:�����DR_����2�������RA�S��\��7��N�CqYTݚ�uB�d�G�hL�!�Z>n�L�GƵ�iЈ�~�/Wf��m?�UO�xn4b�4z#���f�����@�f��ks*����:g�P�Bl���T��(rr��=M���F��F��38:BR�"�L��;��~�� F�M��v�Xʒ���C�錆�zx%���LX�.��\���@%'>���<KAȑbU��҂M���E}�`�����m_��������e?�YLe�:�'7�8�p��"���/����YE�U`�xJ���D�I�ʳ���>w�Q�~\R�0P`>�2C�ǉ�Tä�l6`9y( ��w��A��c����a�f��bJ?[7��48 �3K%!5}�h�f���P7��A8��uR�#4�h�x�H~	��0�d�]	���G�en���ȍ�C���h��L�`��H�� ��~#
vXkQL3S4~�Ϊ�����=�"Q�Z�����>������F�>��F�w�+����~5H�/�s�[�<b�+F�������qf��	���o�K� "�= �@~uuS@ۺn̏��)�J%��p�����ɌR����E�+�3@{�Є�Yne��"yZIp��3њDiq��I%�u�I%�П�{/|�rF��56�I�< ������&X��hw�ۇ�]�,���}ӄ_��tBS��kM�\�;�A�kz�Ո�#�,to��)�� $�s:�К��Hנ�N\l�߻� ��^&$m@^:��r�/6l,#�U��K�c�y��\ �+/�K#��F7�:��W4��}y(.������9 ��c9�����gS��L�B�A-di��3�x���m?e��)F"�C�E�)3S�4J+�<��F�<�e��R�L25�M�e�xb�����X����eG��|k��b�@h���";�w�х���<��}���l��7������9��M�2��>W�u�V��X�8d��1�Yγ�"��d��4�z$�t�u����C�����}$��.�\����;��c�0r������D���_c��)�Qu�?"��?V�P�y���.r�̋�luEN1s:���)0����Q�s�N�a��+�U�x����
��8Xq�M����ڸ-xv�H;gH`n��@�F���0i��5�U��V���7o0� ������=!���:�5g�_Ȕ�*[c���w-�f'�dQB����/�Ī(�%3�vD�,�]B@�5�� f��2bpar��XI��W�H5d�DM�^��z@�9� -�ij������䉻u��I�vDwm��ҟ<[fU��5�I�gIc���Bþ��e����:��RA�����.�H�̦T��5�#����9l��ʑ ��z-3D�(�A����^h�S�h�B�\tE��,u�W��`B&¥U	�I3�AX���Q/�ʵM�����2D�ی_� 9�� ��v�����N(�3#�1n����y���@d|�
����,�v������j����D��~_J�gθ
��ŵ���p�̋:iZ5��Rq��wAq�;�M]��$ﰎ��$�Rt��q;��K����_�Ѭ�&瓋��na����(���x�7��}�U���ic�%%>��$���^�ÆT��E���f�G��.qA��Y�9�t��/<�t��]�6:Degd��8�޻"���%�7�p:ʳm��x2�V��:�����O�^�	;���,�8�����~�w-�	�ޓ�3���G�X�A��cC�F���0��w�X>��T/��ܦ����lAm��r٢hDĪ���6.g1s<5���b�߫ P�N����4ɧ2�ܹn��H
�QK��M�f2�4�����>�P-�Q8ʄz���sn1�ĀE�$�!��9����>��GذB�c��H/���Y��.>�(;O<�z�%�5���P�5H��R��?d��m�Ϭ��#|�0�6}�\�>�An�S�)�͜�HX�F��2�&ݳ
A��R���{hZՐ��,c@�Pdql%B`��&���1�S>;p`i7f�G-9��?,��~�M�\K�x«R�� ^m�������'"B�(�jV�@@�4�H"�-��q�ط��	a�pHՁ����i� GvpXl7#��{��d�e��/�D�y�rÖ�����U�܉�
�G�lGf��<c'�iv܏MCk���w
1��Í�VH(S;��n
�.�Pm���Cb�V�߯�	I�x l�{��;*h�E�v��nE�ң(�Z����J���/	9��l�}�epeQ�f����i��Rmxz�����f��m�I�k�X�+j���E?��\g3�1�M� ����r'0y�t�?F�w������V�jyk->YkX�H�7�����LNh�"��y�$[��t#���̮��A
�)��^�f�W�4TS o^�����k��LU�Ӄ�@C( ��}��6Mxt���	P�r7p��myA�b�fC���:�M����o"M�H�܉�>�/Մ܄o��[�Z!��͙���d�Pi�]Bj6�ޕ�b���u{#�ǌ+?��UL$���y��T�,uL�38��͜�@iM
��q�TҞ�e��+��8�2u��4k�|)�_�tݰ�i~bŮ~j�:��2J&04���#kc*N�[l:�'�w�I~��X\����]�	x$;��=���E�>�r�Np��]:X�*����ۙ���D�"�>3�=,41���G��>�ߞ.<�U#z��:���*%�	-c�l��Wa��?�� �+K��H
�`1V+H�(_TԴ(�M����Mq�t�P>���^�0<G,[�^Mf��r�.���t&���J��9�=\͙��9W5���a�ʚ;ݸ��@h1�e��p4)|r[T�E�c&y0�h��ko��WhLB?�WB>sb���ئU�r�C��]d��R�`�P�ˌU�N���`��S�U�3Ciـ�3"���3%F,;9�~13���G�'k�ց&��\��Bh��e��2�|�����6�6>(jװ��$hT�Su9��(%gA[M�|�@� �-�Z�4z�刻 �M0���  ��+�EU�`Qݐ����i������]VOW���S�����Gٿ�]O�x�]ʾ�ݪ)� �NH�iۛD9	?��l)2�:�.0�u4�h�5��m�E���?�voF7yt�v�����h~�!�-�;nU��m����(0���O9<�Eǟׇ�k�r�e:�f &]�����c;�5���x;U����kW�6p���gSDS�ь���.4��.1!�3=N��e�#��(���-i��t���/}h�h���>DO׀��A+��.Bk�D��N&f:�� R�dGM9��������-��·�U�\��i��Gr�`7	�5N<q݇j�K4����c����c�����ޯ�+�N�HY]&B���t�c�ѫ�/��6���!*vS����c퐢�����K��j���n�֔���{:��Id O�j��W	��˄��xGM�2���R��6�JcSKu)«�\��<�!9~o�s��Q?0�4L��Q	��N���,l�N\��xy�[�,?�>)���� . ?�� ��5���5��r�7�V��p#�ˎ<����e��% c�d��]W�<��:��p)�T���r\~<Ë��bH1;Tg���#���=^!&����y#݁&�������:֧���w�y�o�u}��K��5NrHK��Ѥf���<�'=�8�K���PNj��z�J���&u)�k�:���WW[��Z�8���з�&5*P|L�:k�������@�
��l��~wx�Y��9�s�uX��l�~���r�a�n�U��!��6���'��~Vnr	Zױ�V�*·�{~����L�$��w̱������h���O,��N�`�1I�&��s^�X��`�BK#Z��>\�(�#�u����'�Ɏ�EYE��q��P�A%Ñp{���>oq���(�<��7橠[�l�C�,b�?�lI,���j���M3��ޢڈj%�.��쁔I;��'���Am�~�7�G���-Y�{�'�Cc�m��
{)�yV��m�2I�X��6ʍEM:�XD�
>_��i�f
]��\��[��t���
qХb��<��Ǳ /�]��"�v�#$Ԕ�פч�������.��&�r�C��-3JE.Ë�At^��u
p^�dV|bC梅��U|��}��g?BqQ�H��cAE�N+�;�H�ke���Zb�A}_�[�mN�)�ԞAr���6j��}�~�:���)k4���A��!0:�Iz��`06�
P��֏����±6R�����e�)��X�]�=�S*�M�1��[�a���\boH�[�#X��x�:�f-G��G�p���I����s��_2
�-�B�����4���N��NU%���'���ۼr��;�jkw�&�2I�Q������i-�*�R�NIz���n���;ة�0�eVnv6踥��1���ċxoX�Θ������T��S�0�����WFVk$3�{��y�����tv+=��/vߏ��9�x�`��5{��^�;#	-�௟��������Q��h1)�_���fR=������S���I� �B�2p���~�l�-����.�iv����G6O3�r�����.�,��n.u-� �D��G���+�.�nJ%ާ`?9�y�e�����ޖ�-��nr_��"��:�ֽ�'�ؒ%L�m%���hQO2�ͅ����y5��]?:�Fh�[���SS���`s=����!�����_����.�����s��5�Q5Yg�tl�V���f�2+�!���gqy1�S:��l'�a�n�&.�3�9��������j�G����>��`L��7%��Q�1Y�㑅��݇�>����An[팜
�6'�!=E��d
��7�f����Jf�:��lb��l�,)�'^J�xޝa�V�
l\�Mz�����;�7�w�F�����Jf�w���
WP"�!�����8-?(b?�
��/��T-砀���kM���#�S#�P�Tj�g$s:"X��u^����*��z��ֽ��h�C�w Lx�����puOk�M���|��*<S�O�f\H���b�qv�jM�����D�ˀ:��]�'Ta��dt�\��oY��.
��炅���!�&���SI�`���!wo����Y.}��q*�gWȳ�;&\o���0���a��������*R)��������(��:���Ś���Q����Vʹ96]�y�%7韠v�C+��Ќ�E��s�/��[�T�ۂem4�3j�qV�nQ���պפ�r����Y���t�� �6`:6=̚S@1M�� 6:����N?\����ϒ'��b��:��H�h��
�,S�M��M`�u<fɹtV�<=/����6#z*�;|���2B�d���'�
�h�@c�k3<&�H��F*����ל��	���&m�ђE<�%ߗ���f����N6�̕�oԛ;���k��J��j�R�'/� e_���1�������ա)��ƥ�짍���ݰ8�|q���.��o�o���F�%J�x;M����X<�܏��L��[�ֶ��~��rC��}�Y>C�y�ܻ2cn��=:&9T��g������X�V��P��U�4�����iA���u,?�3������U@�����8��ޤ�I(J��C�zq�K��3!˫���h �r2�k�~�UGG^Ive�"��ӹ���G)�s+���j���z�-)E�QZ����1h 	�B���1v
:|$��ˋ��a���c"�j���؂J���E�~�yX�2f����:<�<H����� ����$�ݍS�]�mBp��'�'���* �~��iq6�MC���-YH���\��_��9e� �(��!��,����%��I���8�#~s�X?�.߇߰�B(��؆V�p0m�]�Ը}���I�ݮ�b��G[{J5�XvЧ�u���^�>�ٸ���h�m��6�!SD��џ�?�Ð셹)�_w�#~X9����q\��٦�-P�t���td7���3���ךf2�al����RO�+gPV���z�����[�H�H�@B�=���b�zrvU���#��{�mL�!}x�l'!�� ҬR*�����" <_�CyEj� W{r�*Ò*J�"�&x��i�@�.j�8�kfI�^���p��)��[*�B @������ʈ�e3���P���&ǐg��Q��� �l�7��05P�T0F�6h�-����{�z���>%��ݟ���p��p�]Ǟ:�o�.����� �`>�����k�e����D�Ĺ�Y�#���8�\�@��Ǽ�1��+�V���YI+P�G���Hm3���*q�#q��Et��ev����	����J8����{�P��3n7Yuc��j:�׽�6�e��3�������B�?ք.8/	`�Cs�V��v���>�ĭ�p)��ގ�e�~]wo�2w̔l�Wvv]�A�$�&J*�l�+U4�|�	��9QL�,�=���<��O��NM��8d&�����ȑ&jbg<[��+mi�'��&��0~�M��
�,1Hp�Ƨ�l��qRt������ȩ�b(ۑ�^�>���SB5\��P�<6�*�;�֌�"wķg��<�`^�.o�/ZT���~�7�/zᔿ/<X�:�{���kO�jƵ����� -^`WoNa=>X�������U�lY�?����9�Yw��=�t	 &s���i��C���c�	��J��h/A����"��1���/�&�]d	�4��iJ�7�� �B2����>���[�]���>j��WKI�2uo ^����h���';Y0G�Ĉ£�VeY���[��u�l�m!l{Yݏ0�~o�Ԥ9��/��j���X�+�R���
���� �_[1�%W��:cz�t�Gs�$ 3Oh�80�nC��uy%����#`f��!�Rql�7����ze�#҆"zе��ހ���n�o�����+vIk�GQ^!�M�O����9�b��pU�#���{��<��^�	@ɨ���(o���` :[j�
h�K�PQ\"d#�F={����\2�Vd0���EǮtZ�ť���	$ �f������^��'�8�6����
C���%��?q��k�~�A�qp>��K�̝tvd#Q�����nu�0-�M���1�N����?�+M�y@�d�2�F����y�כ���J1@��`[����r���<�H��+5I��.uTg�əS$�o�m�)]�O_ n�Kn���e�R��<rfkc�H�gE�}X�oc�%U�޼��/ά�l�Z�*�d�[�qkh�s�J�@�p���5�T+{��a�W��^�i�&�n՝�b�%��m=w��:r����W����D�Y��N�X��_��Z��S��!9�p��Z:���T�kz��	No��@z��})��ܨ��Li*t>/<�lQ~��#�x������l��1��Px�(At����K-�^P�{7�L>Ѝ2o��=�ey*���+MN���P:$v�Id5�'r� -��_rfm}���/�yٹ�(��}���7Qk�/���V�"Q�0
��]��q��5=j��R+�t��"�q��V�l|D���j�M�X,�"�$�>Q�Q���L�f�0n��l9 ��"�����GIS��;����Y�� �?E���8��jA�FԪ�"�5�[F�#����__)s٘W2��gr��)��Gs��Sq�����_6L��n�O4V*�����l�7�Ͽ Q�?��v6
�c��DԎ����-�҈�CA益l�M�ޟy"O�IU��r4kj���6�������v����\�a���v)�(���07�� ����:���ۢ�?���|�.R���E)�c�l�.�]���ZX�I� ���4�;Bk�#Š��>G�}#)B��Cm0�PN>H��R�Ԕr+�tC���X��6��8
4cF�X���Y��=�vn���@�_Ҧ��Ĵ�_{G"E�.���>�	b>�T��?�5��$`e�_��]l�Z� *�@[���_p���.�5j#*��!��#)����H��u׈;�Y���i�N�v}�sH�[���=�%/�{�B��wa�ݛ;�����{)�8�mK	Λ��]�h��?�r����7�,�s$n��H�s���V�P⾼8��!��D��`Rz�6oG���2ۮ4���[P��q�3����#�o8��O�A"PuB��W�V  ���dG�X1�X&���$$[�Rߊ41� �H��d�?�	r�6,O��O��9�ue�E��I$��v�/
,��L�#,�M��=��FE
 4۷����X4��Ԕ6�	}c�ɖ�b�6禀����4!�|V���h����7�
�2׎_0!����p����^#k�Gts�;�DnuMj�Ĕ��Ȇs��`ENܻ%a5��fpCW��f�(�uˡ�2E}g	�yQ�uXa�����v�$��er�|W�_��?�1<�!WR�{
z0�QB�Uv�4�P�.��?�B�'��+n�#��nѡ���|G�Z�p&jRkk1y��0�wV~�{��<=? ���!�m��u��l�a�n���}�;�,D�]˔l\]�>�dr ������($0��q�����?(�@�Y̍�Ja��O%%���3�޺�v,/J����7ֺ�Q��������a��*����]��\�O"�3Eї>�0�]�o$���2#�O���XD��9��𲠎׹�u$��:�0�X���tP�x�'�=R4/W�SD�yFaR�5�����A*b�#j�-Q�aa�
3N%�����g��:��$�V0��k���X����86�
xe�x˟-�Ʀ��B=�5�?�s��	M�DĤ;~��H�%ePD�H���1��ْ����,�Փ���i�tF�*<�"�W0M>syS�I�c������p ��:(�@vh�!��m�Y5�o��žA��Vj�U�Ơ�Hl����j��Y�l��FH���v����٤�4nM5���r^�ެ���T��t��k\Y6T
�7�ʃ5C5d�V�6�7T�zqV-��h�8���$��b��1"̐\/�>?.�{m>N����ק>�=�����<գ�S�#�9;O��zL�7j���b9��l[:�0.���pV8�2\UI��vl:�`�=ǟ�1�/����h�6r����%ŷ�|����DA��+]>�d����f8�`���{���c.���)�_��l��A��)�.�Y;c�RU�D�{�ͪ��i#���8����s��Z���?���vUF�z(�^L��P��
�р����eqΰa�[����u&B����QP���Y�'A�C<��RՒ�0}J��{m@����v�w���"+��<|}.�/���<N~�u��hg�|��oK�t���	�1m���9�Qm��1>t�i����b�r}�6�6�U�3e/oHL
!9���:U�Cj�����hS��l}�l�T*��O��:s�� p�RܿIG	��1�"�R��@�#ybf�@�<�3Q*'8����D�@r� ���茂�ح�,���v�s�/)��k*6�*�1���'kQ���6Q![b�p)�����S����Z�G���="�/�1�y����%�UǄz�n�bM�oX�<1����r�[�t����~@꯵��廳�=���b����S"<�.��ǟGT_��N�	�� <!�JT5�Ur&\(C��p�e�������D�5PkG6��2M�㵏J���L�"J�1���G�q7r�y�s\5���JX�NI�l�M�i�yn\y�U��Tu�PYĲ3���:�{v�LP����!K�"V�7c���,��ѿL�#m�φNW�{
������A�G0Ţ�2��|";&�����uM��^`�`��	G�C�S���o�_����|JR����N8jm:������1_�hc����q��7<_� -/`�V���'n���Pz�w�*Y�Q��F�O�21k�T�.��DI��PL����=k���u�r>�D��[$b���n0�W�Ï����ooS�wTF�I��mt��'|c I�`��2�ϑƫq��y|mT�.���rs_8jJ�G[%��{]Y2r�Bt��p�|���w5nv�D�`�i5Pޛ��f!���M�����S"-�t�����䌽xft<�/����L���r�q[�v�B�q��T�?eҪP���!nr��N�����6+��p�g T��Yz�����A.f�y�3�۪|u ������$�T5ܼs�wP�(�)���ܮvsyO��Z@f�W�+)���`F5�e=�*�wٻ������o8^>/g jnޱٗ��u�_l4�	V�Q:�:�w�����D�5�
o�x�k^
ab�v�����M�v��3��\@q���� M�������u� �,7H&�~<��oQ��ѱ7����?�V�׀�6���Q����.�x���s`BD�Qҏ�k���G�E��a����bӡb��yD��:'��ZȎ��������^r�z;]L7?�8TU0x?�P���R&/�q9y^rIMW5�=��`��0W����S��̓t;{ O� ��"Rh{�<rNO���㔷#��uߝ�5������O�Q�#���󙠰�U��9�T�� P}���_1�<�	�B�%3�H�q��5 T����ν�ȭF�$Ե�q蔷�.���.�U9ԁ�/_�����~�� cǩ�_������P*!����b��f�'I��f��*��[~"�?��db	?����s{�r�,�^����rG^���z��S�(FރګC��p�B���'�V�&?�޳�3��sr���M����#�^�>����+�����,�0�5��7薷f}�?���l�{dn������L�����N�,.�0�Dy{�8����h��Զ6������ �'܂�Ҝ2n}�f��0�-�C���V��g��A��l˝��a�R���/�y�!_$�-��C��y��s4���k��+wRS�r��TrlI�P�����|���2A�,;e��`�NU�*��Ȩ�� �b�F^���*r���T�
�� X/_)���j:�t�SL�=>omS�n�uf5U��&G�n/'�_n��'�#� �K,��!�S\8.��׀'N�����5��걈��3+5=���k���΢��i_SxA�w�+�}ΰ�H��2^�{{��e���TU�_m�{m#�t�n�U)�!`Ƴ��}�z /&�Ub%���ȣF4%����1C�:� �G6��B4���NG���\�s��>L�o��A%Jj�,����u#��{��t-��ϸ��j�.Jy>>�4S�͵��
�RP8�ݺ{�����X�*��?��ȯ?8�7���SM9�P���Eoꋲ�+�^�W�8��/m�����HH�h?f����k�cL;.KN��<��.�� mȇ,�M��y,���G:jL��� 3C�9�5�$���5\�jU������݀�JK���骍�V��$��$M���#ՠ����6��u��R����l49�5�K��̠$aH7�4�g�馭h4;6h߃�Ĵ]��:0�x)�E�U�Mؗc^v����T�c���WUt�ﳭ0����Bu���Y�o'G:%:Md�F�����<w�̎A̹i����R�A��&�Y��/�C�������O�zi7�}h��,
�6�ޝLD�wwj�������dn��g�Z��W+Қ�3�z�kZ�@y2��G$4 ��x�G�����qǲ�o���k��;�0S��b!�1H��a� �8��q(+-�1�X1�fBs�r,Y	�:���M|�׋r�:�E����4�-02j��Ȳ]0�)�_�aި�I��>��:=vM��YY^�Cy�/���6v9I�n�����;���V���9�m��a�o
�.p����!�� e���:�ŉJ��^��![�B�Ƞ�3���2��Gs�݌ݘ�7�ģ}9���@�
_�Σ_G�̴��'� @H(��0^��T�$p/�m	��k]%S���꾪��9U�S�c��3sW��I�)�^Ek ��9�X��d.}xąWMe�ȼ@*_c��(:gH%!N�g��5��X�Ԙ���*)\�5�擢4�߸��&�R˘H��"*�3�ݢ�q�lV�>+�ʈe� �>�������Gh�u*�O�Ө�HyM�ϖ�]��G.���f/�������6h�l�����Ͱ�r��em�qc�"l"�q�2%+U$ÿ�$B��ؽW�ݞ1KQ��R�?Q�@�;k����HcG��
�TM�����(X����e-�̃����9�[�?P&�i��Q������V��������X�K>Ҋ)^�yN!�-ʁ=�۵0��A��O�wLR�b֫�№���A+@��Ήq�:����A�4�3��nse'iQ��"##}�>!����eƈy/�k��ųO.��//S!ؚ��+ߥ��u$ח��9s��i�}�C(�h&5לN�uxr�q)LD]����X��7���������0�Ë`ǌE�iq=�:�Qr�������ep�)�t�/��/��猑�<�N:X�������=��V����OMWI�:p�u��j,:���?�:����u�~�[�\�}��k݌ZP]�`>�` O%*d���잢���Q�}�N�-6�\T�����nq��ZM��]n��I�8$Gsأ3&,h݆�+aal�P�貆���Ou�����������r�Xk�4��^��_R���c'��X	K�.�C����W�A��!�7@[A��ɶ��s���H���~�b�U���2R�>k,l�o.�C$��M�R�p���؂$��M����)���d�~� /R���&x\ċn��ޭ�����s5��a0�yU�hl˙��zg ��~��0k,�̉�5�#�Y�Yz.�"i�⊄`+'E2^JVc)�"����� ԼZ���~��=d���e�:��ay�巧�R����8&�_�$a� 0S��)��f��/��Kbr��>{`EeL�p�R��Ż���*.0<�*�n1�JG���[G邩�+x�1�q��N�:���:��4�	wJ��|���ʯ� ��^Ip{Í��E��8GJ��;�u(A�~y��� ��(0�|��/>�k���l��+ܢ�[�KQ�l/pF��6�K%Du�Q�̷�,�`�	 ��⚹*�u��bxe6?'�j��a���$�KS�g��� G�w9d.}���T̎94Q��'OE�jY<\j���]�)�� �yĻ;3�l`��E��xZ���i��kC�h߆4I<;NWS:�{�4p�}Z�E(��X�-	�ER��?��_�~ �Q͍K^p"*��^:��q����R��-\��]��8��O������� N8���:���5����n���A+��k#L�Z�4~�`���"�L��7�e��6�u+�gݥ[��!ZA���ތ�Cސ|�#`��� <��H�Iʦu+Ӻ�w��A��(
�~�w6���^��K����IĽ�_TQ�!X�Vo]yF�ϑ�9���V�5AĚ���U�=R���йŅ,�Rl`�m6�y=4�x�X��{������X%N%c>B�&׌�4��>��N�l�������*���;s��aM9��[�4�LR��0��i|�V�_�v�<8K%�//y����~]�_[7m�#�>�"�k�<;n��2x���S��^�¦n4�ޛ�ҙ�x����2��]����0���_v��6��2H�W]����1(��`���Z�8�H�Sv}����{��F�{jF.�I��}ƚ���غΩ5f�	g��1�j�M��"��M1.s+n �<���;�)�Hz�3��>��a&�E`$�"6@P`���L&�PUNY�5t��S/���������I�F�O�O�I<�Ubo+��yd	e���'/D����R�9�?�P>�Y��*@u �8 0��&�]��׆�̪�h��A1����?�C�؀�-m�"�d9#=G�v��]z��v�P��'�f���5���8�;�x��,:tAL���oW��a�s�f\Z����h����Q��﮷5�Wsu��������x���6�+^2���4��(�1���a�� |
��\"��ObX���cp�n� �b�a���� �AI��+�}�~s[�}���J��5U��5J���]ȁ�j;��gLc�H�+���H �Ngf<���R��]EF;)�[)��Y.�˞�%��b���I#4��cHӝP7皱-���l����
�eVӅ^��u����r|/Q�Z'G���f�6�y�K��C��C��V�w��!��߅M(����5��\�ͼ>��b�#�m�AY�3Jk;��F)h�2�Oҝ_M�
�.�R峟r���̂��M�5tf�&&�/�i�9�TBbh�:�Vj7�{�8"�˹���u��������a>�O����)(]lJ)�Fp�.��e��/xqd'ε���:t+J �@;dǣ����m�O}幬����L<�}�.?<�k����	�\����o���ZIy��l@/�E��|����9쒡�B�C7ȑm��6�X�����W^� �����t�Z�.BuŝU��o	V,�xF���1����؜��Ĭ	�֎�YX�/!�H�:���f�\bnV�w:�����,�["f��8����?)AjW#R��V"�2��� A�����ٌ����ᓾ�����܍S )$z���U�A�	�R�wey�(C}!%́{�|'Ƶ�{�A(��>���D�Y�^\��Ga*G6j�0�Ӄ���T�=[yd+ACz�*_i̒��d">]#%t�_%��aA5Y2#<����$-�ދ`�y�Zn�A��|E��8�1���jFG,��M^�Ji�.��ó��h7���(�}"i�e��Ў�s�Xt��?b7�g�$�)�"z��A_���<�ɥϕ�� b����\��#��<ۤ:~^��3�v�_��I�D�K��4 S����q	ie`���Ž���W%Ò�K�!��Z����"G�s?�}�_!�	�0������)z����d�tC�~�dC�O$E1�JY�2��A0���=�s̂�L)|��;�����ϞG�t�2rj���|��  y��z�h��[ڊz��ő6
���{9���¨aD"4��?�6�R�(s��Q������P��Հ���|!��	�����4��1ˍ4U8�B�(�: ����q��-��=m�~6Ha�A�{����`�.�/��>|
�:0x���N�@xwE�i#[ri�e-?�[��H��=xOl�!�Z.n��w�(���gH��t�q���-%�Ƀ̨���ӭ� ��b��3gW9Pʃ^���.�r�ɝY%��٬.���S*��s�_P��b���gg����(E���m}���ع���
�,��[��M�!嫦���'�Q�pF�Aԕ�LSh"j�bgp��q#���X��#��(�,�v�u��f�W-���kh\�wT@Z=o����y����������c�&�h94~�R�1�Y���l��ڑ�^��<E�1p�s�ВȟV��`5��5�}�^W�xձ(�c2P��PF������I3��Wctpڦ,��Z���Ɓ� ���Y�P)Y�]���7�P}v�/lg�ÍP4��}[��>��5(*ײPb�"���6O点�]�_yC5hyt%���K�
�q�_#��ʨ��)����>u�	����#qX��>Iͫv�{u眳�*�eƈ�&J�T�{`���}�#a��J��#��ոq9��BDn�0��g8:
�!g˜~w/��NJ����Ψ��9��ɕe��Ӝ�;ҭ�_���Rw��5)L��t$����AN6��ġG��s��]��B<������G�]O�uP׺mR�u3�v��tȄ��G=�A�?vEgZ�F(�{E��O�ʀD�Ňy�߹
h+�)��ĩ 8�.:3|7�64[�k�0�BоL�D��U��� ���6N%餷ԛ�5��"w�$�  �-�G���#�o2SA&���M�S�0�eB�4]u�G���*�aAj������`���@_2η�0~���TY5��;#qQ����4Jf&�s6�����K��U�N�uCn��o?��b(b�I�O�1���\�����;�n^�=�ilAA�*Y�k�G+���S3Y[�*���ˋ(Ɇ���6�y�5�^�A.Ql��K�f9���q���mHC_���ݭ�M{�oIL�����%��殦O	� � -�|,�1�&ue+����[�����m]cI�x��*A�� �a:���s4,Mʖ��O�H|;�� m �<�������,��1��L�8Wr�x_����O�����8�u+�� ���C] <�T��BF#���Eg��ҕ�t"Y��R+��n�u�ymM�9NhQ��~n��d���Jw�7����3�qʮq��b��2�����@�Q"��WZQ2e�-��=����-W��d8�_����pv�q�~���O��oW������J~{b�##uQ9�]��1�BW�tɓ1N�D����y�g-��Q�_*�f0N�,S<�p�����3�H���� >�տ��G�ck0`�h)F:�nN��y[|����/Fz��z(G�X��K�LZ��3r��g�i�jk���'1Q+}�SwD�����J�ʄ2L�D[s��$D�$ ��C���mP~�=����Pc�Q�)3.7�4�Z��'�k�SP�s���ݼ���c��4n�}_��3Đ�� ��z
���tA����CE�l���Yj`P�2�=)������+���_����>������`�����ާ8��֋�J�����ն��p��^�c��qg��)4d��� ;B&�U�Q�����$�G��y����Z&z&�ex��c�6̶�+�+�J�
YA�v����l��`*
��?HI�To�4�7;��F
�?O0��y0'*�;=Kd2�O���4E��0��N���i`<�\K�1Blbյe��6z=ݛ��6[[�����{����Zwk ��K�*��U�_����(�7��v���
�(̈_��D�y�v�xX�o�#Q��m���L�{�I�(P�;,-�
��＠@���C�N!
�+�ȷ?�,e%�J�\��Ж�I�u�6��|��",�<��"v�ƒ�吶��^�E����X�5�04�Ŗɬj�R�j#�ԕ�AA�QT�D��5�ڠ����7\uܩ���L���=sҽ��e��T�|FT�)��r+�M g�@��b��.9$Aw,�T��3S�I����d����TՕ�@���`b�&n1j*X4$�o ,v�.�u������>y`�� �����'p�XxC4��⋲�A?�	�b� �rO踚LY߼���J���M=�����˳������*�:��8�W�M��W>��y�Umᢦ�4��|:gڷ[���3�d����lB��`�Ϛj�c�^��G�I� �v_h�3�/449%�q�Wжb������ �����Wv����X[4�0��7����B`�:~�K�~���<bǢ�.��ƽ���Y�Q��`��a��H��t�������e����vj�����]�l�n�[F�i���t�C!�/.>o����NPA��b0�CIB�]��ڵr]����\�B"�9����j�@h�*����8�^�l_. b�f��T|'f�C������4����ߦ�pM�F�g����)դ�@�����d(c�6[ЌLN�@M�vٌ|%�6U�e��`��Shb�Y��@AD�
ƈN<�I�gb���Q=�z��$����}Rd[��^2������רR�~����ž�*$K3��L�aE��F+��^�T����n>i�=f���GA��o��D ���)�|�(��"���vt+�]l#�}U�A[Z_�$����� �a%�_�X�b�/^�D�st�F��-���_����#��G��8�"i�,?|XE(�DX�@����F��! +D�7Y<tY�X��d|�t�]�g�DR\�I�ث*ꏺ΢H�t�2��A�,�ZUk�����U4m-�ŀ�j0T�=�i"��Z�i�D\<��mɊo9�r����E�C���g���)� ��|ѓڂz��)��v)P��U��p�i��L�b��)i��A,Z��ڧݬ�R=j@�鰘����s�����ת��m�#y7m���tM�1���˼����P(�J�C�L�A����!)�����Ҽx���YތY[��͠c^� �T�E��Z�sԐ�#%.y����W!��\�X���[�KQG2j��m���1K��#q-_v2��I�O_�dҞd��](8܏�>K������pb��w�
��Hq�C�a��~��X�	8�Yݮ4�@tp�:���w�����V��z����������%ó���L2���yU̬k$c&��v�+r[oH���[,'�~���x%S����U�����΃98~�b<жM�P'�<J���ky�w�1�Gg$]/��Əڒ>Hg,�s�M�h�\�p~q�Q����x�
=*����&cm���2'Í��#%�M�DY�Jޑ�)�J26(�� ��3��C�F8���<?����$�/�?{%�S ����,8e�۶G�jvÿ+(ǉA���f��e�~�b�� �<��j�O��A{z�?�}96���ډ:��D���mh���������=�c�JW��~Qb��h��1���_h��e�]��T;�>�Y�p
�K|o�qS��ju˥�������./G�/�(X	̮�*B�=@�tc��ꯀ�Kd�Z;�C4�i�d\�5e��$��b=�5g0o4�I��$�'�ϭ�!>�q5���9dx��{�ŗ\d�ܫ��3h�Wv�F� :y����������N�3����<"�dW��g��b�Db�O��1�}-�+�)�KKE�4����y"�v��>7�ߍ\�}�+���\\��"��D}��/#T��$x�����@�&�H{���esR�6���~ˮM�蚾e�z����9ѡ=/�̞s��;ط��=�n�>�D��������@�\���[�,�sͽ���+(1ǎ.4��bZ��B�c2�p{|���d�жg5��#�\J$��pW9���X���%�5JgV/Ʌ5T�E� <nF�8Bܟ�H����S���D�ޝ��C�U/�O�'�Lq�[(�?*���r0�+�j�߿��$$0���*�� q��� �=�CIOA�+�Eq0�=	��F�K]B��"�n������`�ڲ��ޜ/oI�[�غ� |O K���9�Å�@F>W�����P�`]>��@�h?Ɔ>Y���b83Uy�|>�Z��q:�0٤N���r��j���8o���-��)�Va��>X���ȳEr���<�٤�7��DbO���x��G2�o*�#�W>=2��زs��N��O��>##�2���`����э��i4��5���Ŀ�����o��WӅ�|d:|��'�����'�-Z����,Fw)��S2h���E���x�Ce��Q���|���e�p9�]����q^-j젙7*}�r�Ed�w�)�L�)s��m�fA�3�ʜ��K��EӇ��*^��l�	Oa&ã@z������/����}�N���$;�	%�JY��n28a����93���������=x1,��?�Et�a�L�8mj,�Y3��zțY��?
7Ϫ�F��f'=v��u�͍�<��,�}��|�2l&���@G�����$L�E��F/�Y1BlW�I���؀b��a ��{��S�,@:��֊l��/�6FB��wZ�s{	�����	ʵ:"�y��sI_�^�C�%s�?���p5>�4�$tWw/iC� "�j�u?�k���z,�~�{�L��!��ӆ�I+>^��K���uX�p�#��u`����eؼ��7+�3d�Q\�St�c�Gl?���8 �'��^��Q(n��b
J�x��y� _�(�(���݇����lvx�M�+!<G���'ʉq��6t=c��_��w��h�3����0yO�������в����Jxg����-�F1#"Þ��Q?�@�4��NW�J㯓��ElU��E�N!���knO����ώ|$%��B��������X!8%j���;6�U�i��ܵ�ӫ�n⌎��lnjh}-G]N��R��]˝2���q	p=�_`��P���u� +?��܅a�_�4'���i̓�u�b-hۺY�ѷnB"�c�4
-�������˛Yi�f���v!m{�WU�uE`B#��~[�MsW�w�W��5o��g���go�8�~�J?�V���~���C0� ��|��Y.�����-�
ģR��0ai�m�.�.��2_ډq����1	��$���M�bo�j���f+�+L �)�&�P>J�<���/���`�[���*��JGz�#[��҇�H�/��9���F<ؔ�Pu�4�R�6�|a))uY*����-��."�|�%��Yg�LL�I�8$E���'pS�ƥrq�l�����g9��\D1���ҥ2�g�R�hѪ/`�1�����H���+��0����;*yn���X�$a�Ϯqi�.k�Vx=��i�`��l�K������t&�'R����_��B�{Ǎ�Y��u�a2 ����v1�n�CW�f�[��n��#�@��g�O�go
nk=A�\��ͅ"�x����B��r*��^�2�vykj��x\�|Z�G�E���6]���N�y_�_::<?F
��t��Y��A��H�E��s���p�+�6Rb���q�0Z�+PBF��F �Q��:�K=�pqf�Bs$���2�~�S�*�[F7�g ;���"l�v^g=�񮍳W�2=al���dЃA�c�c?}�L�V��?��b�����2bx�)1a㚤AB�����n�ScF�oF���$�FZ���<^���r��3�"ꓫȐri]�%tΓ���ێ�����ւ2I�e72�<�����R������`��K��R�T�m�Y�'�,v�5��U����ھ?����)�:kT'z�F�!��"�,t�k�g%M㎠bK.�L-��%E�A-�j��X����,;
�`��*ԊR��I���~��4�xˈ�
v��[�BS�X8]�T��uT�-�fT^�4;��l�y�0�sS*V�fH�NQ�EkK�r�4d�O�.�E]Nm�C����u4v�����R��R}sVXM��	�q���y�~�X��fq�a<l��F�)`��ɥ?��J�H�����c0��zW�Y�M텱���"Yh�� Ʃ]�a:��X��a"¡NJ��̝i֧���O�U�ZģV�y��".���ẑU$~3���uL6�%��s#~�6G�-�`4�tq�0�U�xr�S�x���3��)���#�� p��̶�r��zK^ׂ�S�bV���LK�W�U�٠E�@o��B?�hJȜ83��#�\�lh9e ���٨�S�ۯj���_{ @J,���C��I���
�^`]HS���Ȇ��`�7�=�.3�����N�'��b�a_�X��z�����'��bX�T�����l���{t��ȸ������ �a8��ĭ�k��u ���hw�)���+�l�����1�����?��fC,�5{1�@T_m�:�(�ky�e���>�74��u�UQ�?����)G�7�a�/���kKs/�n�*j�|aE��TX�9z�e�ˀ9��-�����oY�d�~�&����@�f�R.=o�^�F�Lt�� vD� ��`����A!�^r�qF��cf�9/�Ey��x��-xJ�P�I��D���:�FlG�~凚�GP� Ż�� k��__+�15 ���x*�3�|��C�@2�{����uǑː:BǂEu��K�AIM_���Ji�B✩����9��KL6L-8���7mu�5�d�8�UzY�1�ﶻ���hѫ�� ��������X�~�p^שS`G�UD�.mA��K;�B�]fVXy㪭Ut1�w���+��:1�L���='��`?������&��Ʈ��WN���3Ep�\��B�LGH�pU�6/?��.K���;	���fu#k
��4��0`�YPx�����CC�������_u��	6~�"O����r���l�#�[���i*Z|��� ���Q�?�f�ȿ/=,- ��*A�O UjN~W[sA����4{�8��&!VM0���bm�(�y6���p[%�3K$�_������Q��|�6����t��hni�N��N��P�&��WΠ�>{ǆ����3kOX��w"��y�E�S�!�!�9��� c�,ql+`=����43�G�h���p-v��U�Ѐ%�S������d����\���~az�Cn&|y\5B>�e����g��r��5�4�D���Kf*6@7����o�;Y�h�8��C�YT+���f�/v���j]b�5����{���T��q[�ᳩ�?��F��䵮��ѥ���þ%"������x�d@�h��	PJE��@��/g�m�59CL9�6�J�`�n���,h|�Zc��JI��*]��*�&� qXH,��m�2;(ot����է JJa։9��zS����@�0a�~��a�M�Gn;V����,���#u�fK��bK�ڒ9[֟G�������R(�d�ͼԕ1h�),)�B�d+D���`͓���l�v%\�����-�[�I\�@���Ĭ^^<���D��� NP���"LFv�>ѧ�v���z����E�A]_O\y�[���(�ij���e�4�~�m�C���UYk�ǈ��u��^0>�����Ο�*�W�@O�f����@�� ^KȳDǂ�ݓx\�Zk�tu����[���A��K��I�b{�o����m�v�i}�Z��>?��հ��-)�;-�� ��Vv����ئ&eTOIf9�$��ę���BjԈd�i�}��c��̀��S�Y�E	����[�YY�԰��_L�A���nڟH��1-����U�D���0PM�_��paq�W���#��+�D�5)�fD�^jE7O*�F%�iw��>���&?Hf#qwg��Z^��v�6Q�O��	�Z��Ul����d]�tN���%�4	�f5���Wڒq�R�K���9!�xCy�.
I�M�uR�	��;�+Z �s����NX}�ӫ���v�>���ʿr��F7�M��K�\@�yb�T�jwҰ����Q��
�X>C�;���ʧј��X�2ea�Z���hb���F�V�0N0w���Pw���)���X>�2�B&�\d��R�-�(��0���kx��h"<z;�'�L��uߴn.({6/��4��^�O %�2x��i�2�J���N�S��?���},˲�lIn܏n׆��ܷ�G�i~��Bp�3wiM�A�+1�������|��5[I�f��-m�\�n�|L�F�٘����$�J(�	%^�_��w��?6u�kjx�R�b3�f��
�x�d�t^,x&?�m�D�)��(�~�0!^Ӷ�V��L�~�ף$��]rʡHX��#�5�S�(���^������cX��Y)z>UG��.S�H���I}H�&�OǷ�����J�T�g�S
*�.��9��/4��,�R�g��K@�t�MS����N�r?��F�c$*��p�v��0�~h�aT6�8���
/-�ԝ�Փ�dAVع[@6�uqIĹ��B�/��Qp'U2 �*��9��v/����V�-�?�<ߙB�4�s���D��0jy==������n)XsQ7U%K��<�'@��Vļ�O��nRe�-�Rh�o.�������n�ϙ�Yt�8乪\�P�6D�E��i4/��v<<�l����J���N�=J�8�������h6)y��J]'��"�
k�
�E�s����=4�}z���>������FV�|����t�z���+�����̀��Z8�^N�i'+�)���g�G�9�{������ x�\+�H�8�ڑ�x18��$ظ˩JY�����E��9�;��:���)2��u��3��L�����a�=(2ݰ"��E9��˛#�!vO�п� ��<�5��g���=�T�%b��fr	Z*1�x��q�Ȑ��>�O0�H�P�����~F	=��|�2�����f�ڛ��A�B�7 ��g�J��U{yd��g�Hݞ	�?�Btj"�m�R�ƪ��N���ƻ���ʖ��HqɈ;�0�!�7&^���վH�~;D�
�E�G�r���?I��?��wַo&p-���cy<U�R�o�䮑�x!ĝ|ԙJ�A1��9��*��h�^6�?d���L�^��@iD���D�%�w��W�J~�j�g �������0Nye� y[^��<�^�0�e���{��m4jL�Ô�"�_hI2D����3�}���Ư=s�%���@�����v8p��h}�,��5�fRDA��4�2���-<��#?[A��T�͊�Ζ��W֋twJ��$tG�9��6�6�@��>����~��gX����(����<����5��+�(��g7��9�Ύr��#��h�]����x$�)�FY.@�����e�r��5�`Vh� a_/*�8!�4bƝ����J����D%K�L�̘��FR��ţ�(.Wu�S��D�b�bJ��61���b�>��܋���0�=TKO�/a�nl>�J�i�
n�^9^�k�UTR����'f���#������cR<�;�� |6�V��Dp��C� D2U�_<B�t�i'�U�+��D�:�4��upͺ̓�R������Śf��"`ɰ�B�k�d��4ёv  T��Z�TX�Գ��s�g����e�iCM7���u�xމT�DZ����͖�y�"!n�O�$�S����T���V'3yh�_	ٖ��&�nY�,m��f�Q?��;��u.-)^V���n�eh]r��J��h]�~��M�-��/o.%��Aд�T]ʻ2�[���;�2m^|x��*[�lY%�zP��!Ψm�J��H��i�*2���Y�xef�Y=3�[#��װ2�a��DhdP�'j� �55,�S8��A�x��щZ��F��AC�H�%Vw�$OH�|q�Q�8c��Kx��$��8���%�x���VrlE=��L׷Y*U� X� R�,�s,�|aj��o���������L����S�hS�L����k*%Jw��0'e�y�F61L�aF�l�|0lЦ8
ج��Um��lhƫ��~�]�$�x���6�c���J�*k�4�G�M2�ջd�:/U\M̟���޼&"�ތ�n㤮;�O���3�1���Zy�ċ�nģo����\(g���e�G�9Dt(mK�K��/���'����O3���ǘ6n+������_����+���ه��:a�7�Y��t�#�fC+�iq���������@D������V��A��2�ި�C/_�$򈾎��L:@��=@%)&�!Og��є��h'4�`�mƣw�w@��H�s��+(˱A���;	���1x��_w�x�84�{/O0�t�wa����)��]������B�>졟c�EgA*/���`����M��w�ֳ�RE�,�3Yb�
�/i���}$��gQ�ܟ�NB�@<�����K���/���3����c)��i���c�qMk�70:]8y�jL{���}S��z�#~��f��!"��Cd1j����LCҤ��$U��w��S`#�,�c��FM$ ]	U��D~�hkcذo( ���+^���Ŗ^���4�"���J�Af��c�l��u�����z1g���?�1d-!�t�]�8����W��ʷ�wVS6'�����[鼫�$u���;�̂�QTe�,��p��m�_aCמ.Y�!XbۮL/������md�25�퐛��1��)p���c��hHU���ք��� B��M�_zn�1\���-��
��
�h��'_
vm���G��.Η��f�m.���˫
�J*�,��H�3�v�b�m�X����%�<��E��ĉ'�[��uϘ^k!�c�)���sg�&�Cg{6ܒ�_E�.�V}f9�7�i�\vH�Wq�R�p5;$�+9,���/;m�LZꂣ*����U�d�w^�L��T�s�=}4���G�Ҭ;�]�8u�Dv�F	�%����jO��\��VB�=>�ik��V��[6A�xəy�PN񮃢*֝?=ώ���1����	��E��<�o�����.T��i����>����@��Yw�g\D����ÂI�+�+j�]�6zu�Q�����h�3o�<�D��N����o�#�[s�Gm����������6-��|����A_�~X3�:� �\N�p��p�������A`��^B��;}a�n�=.h
���e)K~+�'ıq��D�.=��ک��: �P�ݼ&��Xy*s�rrR?���~ ���Wt�(o�~)�QY6|T(�`��G�s��ۦ�絙�c�C�Çc���wqfG>A�>v��'����J�d�=�B�`<�����2Rئ(�����P�����đ�#�v��I��S����*8��CC��R�޵ܯP	_�
�$��!H�c�./��1ti�(!J�Mދv8D\��`}Bn��F	r<ˮ�������ƮeD!dp�P��j�.�I�s�h.t���$��%�9��J�؝I.��6;���S��������礆� 0�ks�mNG9�\�A�+�f���s옶�|w��[�M�?�qM��}�U�IE �?�p�qw9��E�ω4
��O5}F�JJ�J���&;Q�ͤ�[8Ł`��ŭ�A�6��Lb٪�>�f)�I�����FOn�k; ������9c������ H�8���0����6X���*J1�9����|��=ݨ=pV�����s�Eڍ׮�l��t�ì3Y8��8ڄ�E��ǒZ��!�C`�`�RNeW�SQ���5lh�gzo�Jjk UxE?���5��vZ嗤��ǫ�j���	�����$xf�;��N��h@����YO���C�B&m��J�K��շ�"	�MD!N����foG �?!�\�[�JK1�lyu�;�Y�Wǳ�U'A�S�-O�R�6���m��4C�o΋x����K��@
6�p�9ra���A��Xn}���o��-�����Q�g|L��W�Y�[�
v ����EDk`	�Sba��R,
,"jD/)��Y�&=�����s�vS+�w��)L�y�׌J��'���K3�Y�a�Q�E�.xX��W8M�������kK�V��Y�ȅז
ݵ��=q=Ȼ��;㔥u��e�-y�ˋ�$9w�[��� �^�	���K-Q����ي`U��ލ3�������m��(��D
�L$F �R_�����9�DZ��2%��KtH�j7�z���kt"���^��6�N�ĩV�i���c��Jr ���oцx�V|3��K�ɐ%ګ9�
^Fa���v�@N8k]�S�P=�x�V��9]�5��
m|�Y�'��b!��)������l���*�����WԤ�Ǽh���ϐޖ0��pc��PSo/B�h�`�^9���'?��jf�aD����7�4��n	�Z櫿 �=�?TRY��di¸iR%!��^����U�j�-�Sc}7�o�y��lQ'�s�,=ߑykV�h�� ګ�[<Ǵ�\=M�~mmv�<��Y�ڵ+ǲ��X��p�ea8�7�+���gl���va���o�{w��Rudi]zO��>l��=�K12��!��_��h����O�;�C�J˧5��2 ۖMԳ?eg��A��g���ù�:\�]��"��G����N�_���:�]	C���}Z���+�����G4��@�"Lkgf��8�9�۸�@g�'��Q�(�y�M��p]�lP-�x���[e�z�w�0��.7�}o�5�'y��v�s�f�fd���������wW`������c'��0��sh��=�(ilC��,SC� �2�$^�{��|g	W�@t\�ޣ�S^����{E�Ktw)�_�V $��麭��*e��W7ܾ2��Zʧ ��qDTN�D���X���Q���zөhE-���jYB�=z�6tr�r��W�mR���χ1"U�`��cx�_�
nTI�|�w�럹.4�y�``�Yy�Y�����@�����nSǴEn��(c<�h�X�\/�T���>Cc��;"=v�/�g� ������g�p{+'_�Н1�m�|
t�K�Rb�[Pq��v�l���,�m��8�Ɣ�:�V"|����ֲ6]�e-5�7���eY!Ciy��(M%V�w9).��u�(k�KW��H?l�D��UAGXQ ��-?��mI%������ ��q�Z�����`��\F���h���OՄ�yau�aG�뚵���&���Q���5_�:��%;r����K��������A���H�dfVzߓ(H�WḪ+B�������B~Toِ}#�r�]'!����y�B��fJ?�?�*��ڲ�.����iXDo;͵���L �3��ސ����L�9NVk��f�25�,h��ne�ǫ,֩g��I.b�Vˀ.�R
���uur8e-�cM�WZEԤ�X �2��&���S�y�=4� JN#<�.Yq�l��c��+�`ƻт�kLX�7E��ʐ�ߑB��bD�<ECH��J���$�dG:a5l��\8>��Ϸ��,��&���'�3A!�t+!��H�F����<�%ބ��T�#�G{��?��L����X5�/O�������L��$����L���xP���촛�ua��[�2�@$��Q������!���z@��ݟ�&_���]�&��>C���vM���|0}��2״�թ���J��?R� #��X>ˈΓ���#;R��i��5(v&��bݝʌas�#�0��?݌Ov�	\8
�jB]���=B�����v������jp�x,�%o�7ESw�.���t,>v��b%�}��+عuv'��9�}�z��!aҜ����^>�3��x&P20@<�4��f'J�? �]�Au6��i��YﲘN�ܖ$��=L��GC��}������f@�lr�^�^�^�r�KB���G�U�߿�	���iJ]x��"E�K�Nz<�������zs�w�>��6ת���gt��d8�:��k�[K������n������� �� b9�$�i-�M���p�>pH��Iè|��;�>�E��^*	u{���n��9�>�ۅ˝v�C q��ɝZ�gZ�n��Fty2���A�����O�����P�fuE���H�9�J5�Ny�Y%��MS>��L��^��Ly7]��i���qy�Է1�+�bT#�Ҹ�.b�������{��j���t�3d)C��!'�4/I��
�l<�BMt��#�����NѮ��,��$�mlN����mF���͵s���F��� �F-�<�xI����Ƕ�X�!��jc�6��E-��EM��c ��S�G�/U��j�;<hK�I/�v�C�mz�N,���i����p}1���xecG����-R��\�>t�JU,cݴ��AE,o�h�D^��J�X���I1h;�$-�!@^W��M�ŋ���@n��8v,�:/�Z��FӁ��q]v j��b�O�#b�f�7"nQ�T43�ѷjc0�M�ڴ#/����p�ϕ�bw'�tAz2�Ui��ݫ�L���Π�>73ut��"�:?�d���U]��v�қ{����}�G�
�{�p&�fs��[�]�6�Xi�h!B����|1/�
'a湅��'��Mu`3�)�v�ޔ.>܉.��V1��\�`q� 7�W��.y-�v@�熼|�1I.���R�8Qo�����������u{,o�+P'����ʩ����8�ï�Y��<J�ŋ�ہ�Y-�y�������M "�N�i	�x��|����?. !���'�+N�`p��e�R���s<����t���J'A�+�UGJ�Q;%��U˴�L�Z7�I*4S,���o�"�}��
�xp�ad���A��E|�o�a�K�C����՛i/\x�o��d��@����Ȃ��Y�ʩJp�|4ݳ�aB�y<O�o�ml�2�%����V���X�)��i��~��~�N�W!(DX�v�yO��D�U#K�-��W�9a& �<��� j��.x!g��j�׉I7��PYj�B2!L�D�7;/
���~�����c d��K���/u��|���%����ё;$�i��>v#ȯ.M���l)�ї�4���U^��F����[��|���;��=�^p����j睯O2�{�:\�)�۝�#�Q۸R�+����u�h.ړxw 5%������4�b���ԘK�`��V�Ti���o'� +=T��ui�y��ց��d�S������{��J$�X��{bM��\,�:O-�'�vۻ*���'T7�\�OW\����P����·����B����
��8.�5��J�by�[�������*?�+OZ���c��C�����xy�:�)���Xʖ~@�t�7X�۹Q� �C�t?!����h�2��P�-$���rb��n�"	B2!�M U�ʇG�-Ţ*���w�/Ю�����K���j4֪BGT�L�put������O��0���B�Q���c
�|��H�mg{�]����7���V�ݎu5f��c��x�|���� �m��T�g�.�q+N�'Z9u�" � ʹjk�ho����$�3�Č�5�N֦�����x�?��,3��eT���9ʥ�5YIm��x.3��=^�ʗ��<4x���ac�"{fB����n�݂+�t�'g)���aɲk�@�$XRA�R�S/��&�6�.`@Balb�	D�b�^Y3�:�O�AB5Nq"_�6�����~ˢ���5y�W�֝�e���#�d�
q�*|� GT��y���ż�6ZNypQ��·�9z2�{��<B�R���#��N]]�雎�u#&�21~���uj�%�������wԽ�~Яi���l�q����m���T	BGl{ �=�/'�d��7�PUH����E_q� 9�yU�|.�Z���av޷F�pcZ�a��z�����@��z� ��'�3b*~Z�U������#l�����Z�1�1Q�X����#@�,,�4n}�s�؇-2�&�T��Tc��זp�۰�l�^g1��4�l��������k�h���
�����8n�-E��_'�T�d�z9�z�([ NA����!�$�n� ��U>�����7���%]�}խ�q{H���}gU�,%�LY<�&�����xwDpSL"IPo��#�fS�h�6��⻵E_OB�-*���_y_)�<�j�AeEmn��˜�~������p΅O��)Eʳ�C�-�h�a��!����Mi7�&Ȣ�,=��W݆l��ZZ$)���@�R�����(�$|��E����IOB)�2��ۉ!۽r��x��b�md�l��ۿ���>��>Ć�>�4�� ��r�k����[�U�G�+U�E��J��+::�X�z18N��� C0S /��	Au�ԙ8��Pt)�K�8eK�ѽMD�88l]Ի�K�SMDd�.Fc��'X���]@X�FY�pwT���(�q@�n�MZ
�נ$|gJ(1�����a�u/}��x�S��g���z��g�o�����v:c���2W �`�Q�Jd�Z�p��ި|�ّG#�A��eW]+�,�9��N�D�����d�C\r'	��}��������Z�o�h#�ab1Sو�Z�"c�BM��b�B��.��S�?0U��~G$\��l�w��	�gD78p)GM<c �=����{.�VM̳��cV F4o���?�n��3??2�x���!�Bx`S��C����"�]�T"v�:��(G�W��m���e�C��ݗ[��]E���f�*�g�`��jt�*ѿL��9Y���"�`n�i�u������c���m��vb���!������ǆ� W�P�=}qͯ�QV� ��|ր�cm�
����:�Hhb��R������#�Q���=�JzXF�S�&�%�;� tn^����ڃ�	�:�'���,��)��ϟ�C�ޞ��y�O�PD��y�;�װ�]=ZWn��)X���2�:��Dz�� ���N�T�6��Dx��W4}1�MiHc£ə1\Z�2�`��4��p�Awuk9�W~�~�����$�ͮ��HgA�D�|9w��	]��uDkw����"�b�>���E��:��]���� �7��V(�AK-�n^�͕�RS� O`��DV���k��Ӓm|�s�o�A����1��M�&X��!e�@ՠ��e��3yd��r�����TX���F�}u�*�&��1�f�-PR��08��znݒ���CK�j�1X]�cG��B����;w�'p�{5-��Ǽ���M@��H8���g=���MȩV��[
K�8ѧ7��Qr<F��3:Nֱ��&�y�'�]EtD�\�s1+z_E��qd5�c�&�+�?�&179�������č,Մ�It������zQ��J�R�W��j9ڻ#���P
sR?r**�sPIFVB�:�u�]�Z~����������Rt�Ź�9	8��h�<%A��22�fJ2�R�B�n����ܲ 2��U&��h�#prq\�e+�zr����Hu"���,�#��	�Bw�`���i�׮O)�b��>������Ļ$�nG����7E�>�ig�w͖�"�1�.3&�ɹM�)����zao��x��U.52���l���A�0aP�V�{���W�����&q�:�'����Lu�bu"p����2-��U�!�*���\7���$����8\�v��S��$�����Q�"ߑ��8T2�W�2-���#���,�v6������C�� �|��ƪ"9$Zb��x4 	�k[R�&_�h�����%~
t{�LX�>���T�#v1���y�G�El�#w
�v���9������K�J��w��F����(ÓBw\ �<J������QH�.��7��r�Cm�fi"Vi���,�i��2ٽqA$�F����lb�p�J�R�X|�m$H4UM%o�IW��� 討K���~��ܙ�g��ߕ��pҼ8�^�|W�=Ǖi��!2l\�y�l_Ysl"�R���ѷ:�H5��}`�&R/[��'��~Pm�����v�,W�s#-���W��<0&��eyNw��H����.�nC�#�	�S���REb1�dY�������Z(�h���󎈒�eT��:�p��fas��ٜ%v���	uGS�KYM��K�]�c��C���I���Z�4>��|�Y��#U4�fݡ�ь��w�3��/j_�'���?�v^k�1Y1H_�u!����U�������x�G0�Ve&���UN��kL��;��l3G¨��@��3�N�W�58��s�o��J:�9W�����Jul� ��2s�}����u�$Xb����wh�Qq��g�KOt�x�#����Rc�dޡ��>�{���)S�}}�4t�ٮ<�.�n�}�TG����0PV���'�9�&�i6�
̊Y���CUA�I0(Wc�`����8$t���pt��[̰�C�M�j��� ��\�]w��	Җ���,|pWQz~�1V�cw�Y> ��b��QF��/ɱ8��4�v��W�mo����C&�i�ű��n@ܭ��/j�'�YA��/b�Y!�H�Т'��t��"�f��wH;hF ,���'X��vL�A_��ǯ�(V��S��R���&6WS����@p01	�'�����\��浧66m�&�����v�H7��d��]���-�.�l��0��+�C)Z��m�J$Y��8���_5�R��SFŢz�^Uȩ0_���	Ы���?�L�݊m�( �84�f��`�M�ih��H��n�l�v{J&�ֈK��R4
f/�ašX��鍶�/=��ܛ��u<��~8�a�//35��ǸQ;O��2юUȎ*c�u�haU��w�iWz%N��_;� uʏυ�7}N� &S�|�qU���̠�5)�r�i� ��b�1����ݴ5}L�T�<ҧ�5Ш���5�{��&��G����ԇ�+�O�w�j���H�w�P�{M�R����Uk���D�������A���3i���d�ݩjZf-p�u�;�)����r��]�'�<D4!'�	�WTi޾S��7k:�i����W		� p�k�.k�k����[f�7�Z�h��;�}^���J�(q�l��(�ǃ5�w�C)7���h�ߗ��Z�P�����QJͅM�-Ѵ�V6k���?뇠ם�vhl����]��ؐǼ}�G�G�$�Ƚ�Rn��H ��~sٓ�ɞ�4趽���IO@�{H�9�?S�<�t�T�7���L�3��p��&�c˜�>y�=�^u�"����wi�����M�Ά��y�m��w�6�W_���ruxW��\�sF�z"��h����^	�j;��mD%a-(����Qn@:�3D�:����H��\k?*^Z�^Y2���xjD��7Jw 
��@�;vƅ^�$��+��Z�����iU1�kD/Rke�,e� ���岚I�.of���۲��n�R�w}F�t�0����ط�|i�!�_��8�%sȭ�%DQ�2��3i��1�Qn�"��@4<�#���,Q������$�G=�[�P=��D����3�j�c��IE��vuRO͂I%}G����^�����*����,Mcp7�/��'�'�ŚJZ?z�J�\r9�^��� )G#����X?������֭��暽�av����t��ɭo��ކ�G��jX^B�w�����\�>��?Y�/v���=�'pQق�D��n4�
n�6Nl{���s�u��eA�w�z����	�bpA������K�;,�o	
���~�� ��KNZ
}��0k�/�7��G=n3v-���T,G��O}������e�M[����u��1�LN|��gӢ�1���}����'���-^|�֔CWj�Fe5���740\�!�+��)��|"EߔjT,�n)ʷ4��'�iR�<�>
͖i���^Խ[�ӸX@�1o��FB=�5���{t�&���d|x�����-�U��
%�/Ы)Lm�W�f����"2�N<�J�Y��k��[Q���e0N>p>�ƴ�I��T����>���2+�,::�D��2�O�۵,�A�+x<=��s��Tp�^(�)z�ߍ+��wVץ�L��V���G0H�y �"� 0���9�o.b���&����=)�K��,]V�FF�tc������熠��]H�oy�]�}�ke��k�UF�p��E�&.I���;�$<�'*YOz�[$�����b��zB�+[}^��搦d��D5�'�8"6D��~�t�$砘�p0���;E����:�k���T�MQn*�����G5��42ٗ�˜C&��-3�㚌��{~�u�bx"%����T�ȳ�q�)i��_�� Sn��L����6.�d�5�Ƭ�6��TZ��CF�q���Y�r���>������ė��a@H&	˼b��Ē$��q��h�>����r����8u.q���e���z��2�]�R[���i����>�9��^= ��d(�m�i,:)
������v(4L$I��(˛�dl�4�j�u� �i���P���ȭ���·x�R��\
�ygP.�Yt�V*
"d���u��~�T��4�M�y�4�ta1"�q3���Y������@�Ov�r�j�x��
�J�7�q)��3S�V�� R]�{Wi�@%�4tcA�Ƒd}�nhz(�I9%���7"�J0㡪�U�����g�>G*����$����l�^m�@���z�U��	�<:�����Hc�Ē}�.I�Jަ)g�F�2���pk�aej��闊x�37f�����k�I�$x���e^H������'���\Շ�L�o��F <V�}�̮�� t�n�D��tI¢$���´�O>��ݻ�:�,�6�b�]�x���>��}�?�ݦ_����䆪�7��J� ���rB�Ho�Q|��������Y�����Ҫ��XZ���K��\v�`��F7.��6`��0���$9���3��Ͳ��2/�{�8[ک0Yk���nl
	���LF����q�O�[K�m�!��RϬ1�fi�^	y� ʬ.��1��h��W9]�Czo�V��L��e��u�e*^BW�"���Vz����(�Hu\���v��X]�6��,��7t����w0�t״J�E�n.�my���C�%;���
[��tiv���ŇQ?qv��ʋ���7�ө��U�<���?�pnE��i���ޱ�0�V ��$�7<>o�� -[�R��\�0�֎j��*ӯF(]������m�{Q4� �̆�� o��*���L�:6����27c�I40qDS����+n�K ���0��n0��4���ǂZZ�%�D|��d,2Oװ����Y-m�yH�����7�7PfR�vY�"���?e]cG���Dl�RYE]:���N����Π/s�=u�-X��'#~޶���P1:���;�aɍD,C���R�H���j�I��S�«f��V�/R9�3=z�BglZS��Aa�s`���H8�n�H�����-=��3
U�:<����.]�=9�3��Lֹ��}���l�Y3X�"���	�Ɲ�$�z��Lx�d�"r<���^�6��)��?I�K�B�%K2��ۑF`�q���1��;z�i��Nb *ǝ�R�MpQmX��^ 73�' =0�j,�E��?�:!�d���Lu���A�6pBeEk��ǁ�k(���)�+	w4�eI�6�Pcj���9�� e�@�T��z�%\�dF�;|P�2zq-�sLh�;���&�bSፉ�GV2�/���w#Hˍ#�6������ ����eS^^��[w�-8����s��gkג(a�DO4p{�Q�{�N@������V������ZwhB�j���-�:����'������gY@���Tc�5~QGb� !�_��/��m=Ͻ֌�!�E�����ZGMZ>��Z���0`���hd(Ȝ���Bu�lÕ�H����<|��^A0I��"�p�H�)���>x��A]�r/IZ�}��O0�J�9�4���Q�*��9ɭ��o2�
X��yaw*��I��j��)�
S/H����E��w	{{�9X�+ڟ\�¨�S������'�|*$��u����;�S��d��t��Ll/Ds)�E�g�&VG��-C�{5\�x��I������%B@����/uI՞�؊eA���rb����{l�N��w.ą6�c%��n?����U
��I��b�H��W|��jG�_T^Z��m1E3	a95��ɸ��s-��d���y�Y�/V*f�B|�+˼o�E�Ȩ�lw̗�8L��x���Y��^��#y,[�*+��{/�П�b��r���Ҳ�����nK<�I5��Mg�1l���c/,p�̴�em�@'�����O����<�9�.���`1Q���N�F���@:Q��E�&L� �A�b?v��Y������(������B"I����q�I���#I#��z �Aj���I�03�R����(�Otݒ�<,ʉ�Ո�@!�[�&�(%�-
-s�
K�����]��i��{Q�a�/�Q=��r[բnjѮ��vੳ>g�Lf���q�f����� �d���h��g�f�r){}eŨ���r��� υ�ٔ&:���G�ǳDӐ��p���E�K0f�E��CKL�c�/�m�Rg��Z]^���[z2��'3�����ty5��3�:���)���Y�V�fW����D���}Qϧfz<��D=oT[�n�������H3&LV�9����	�W�fї,x
|we�"���ɚ���w��`�.8	�4_@;�,�C�����1�7�#�3�i7cf���b�vd��К|T �l̻,�k���n����I|[(]�B�G3�J����6�0��?aCnw�$Tj�RQ쓶`�k��`��0�u�����O����N7�t�}���L�r�'�j���M''���������|�Czag��S�t�����sB� \�x0k�;�&����y��8j��Qh���Y�� ��m(L/x�U��_�<��-KI��r#���~ł��V[nT�G����޻�(F	�R{�W����O'ie�WCy&"9��^�A.�H�,}��)c�S�Y���+VuL'zZ���P�>>�? li`y�O��Kz�EE8��a���O-��`Z<�NY���*����,��	��M搣`�0�)�^שEvN�(���!�te"�Mm���^��b[
�]�`c�*�"0�fn�жHj���-�`�~'�	2�-\E���׍�w�Z�2U�T�
��5�nZp������5jZ�n�}�����`�TZ�!$�u���&7��*cz�2^��:Wى�aY�C���ۃX���-U���&8w�$3f���bW\.}�l�r�b�5���D��4�KW*ߞm`�e��aq��݄ZkN�=��q�o�E}k�sq���8��"��騽�~5���iIҹ�s�$�m��E-�&5�d�ܡ-�B|��A��XaS��6����5eqӞJ���ɖ�L�r̷�:�
$���u��@�����)�4���_�/Js�>�/ME2��,��1���� ��[9���\B�# s��$Lמ"�� w��\�Ab��v�#��W�/�ҁE�nxaӲ٣��J"\�^ ����\��a�L�� u6�����G�tԱo�u(沠Ftv�8eI}�V�\H�{�����~��#�8;5c_fi���ɮ�b>�PeVil��˶	����p	ǟba��I16Z^OR�'Z>D�*���@X-�����w�I'����A�&���a+_9?QGsZ����T��C�q'
R˛q�W�0w�LtBK��\�ULM��p!�bI���o|p��-�6ܳ*a$�_�=�À����U��6��c�s[�q�@����.ԝą�`/��ck1Α'=���W�rX� BFc��a��%���7�jg}��V�..���ڇ}��
,`�yn���i��#�ښ#l;qg�x^#���@���3�p�y�u�|6*n�����
ךP`S:�s��nHe�^��.(2������k�T3~E�ųת�y/��A��a�S��x�Fgy�5�=(p��=���"����C�d0�T��m��Y������e�s[ؿ8�(@K�x<3:��$�I|C�x�RD�#�\��=~�m� f�BÅ���%Ό����]e 1tJ�^��#���Ȥ�`G��hD��k�:��cX���e��}Rv�ѥp��P1^��"���h�U�P���d�U|������K�N
��2�A�A�͠��"�a�"P�v�B���r5��LR�i<�M���^
���Qx��;��7�zu������@EYjtb$��Dl-?�<��]��6��w���Ixy�'���MM��9|��I��^Z���br����R{2'컝�v���ރ��mJ�;ۭ�=ӻ>��Q��ѭ;.�gM/�]q��o?Y���I6���e��k{[�wr�'�d�_�^�n�Y[aT��`��|�f�b�>x�Y���,[��r@W��hWd�� �z����O� �e_F��O���t��U�\e(�� �[�'�~�$����ˣ��?��zkp	�UNZ/L<�s��4�'���K�����pw���ۭN 	'4�$y����N�d�����!,`(�w�W���?�<v`��%�ޓ k�!i�"Z�>EfGTmBl�����hZ=��B6���ZG/X@,,�74�69�����<Z���m��0������Ų����v����Q���'5�l����R�`�
���!>=��쵽KZc/{��=Q�i� E�͍kD'��6TL?9��5������+�^GӚ~� S����7Yo�2-B���gY0�b�5���Z��$]H=3	�&�VCg�ťB$� }�m�j�J�	��܍�2~���NP���R���4��WH-���>�B��.�k��e����n���N��"��/Y��pp$��ݘ�a�	O`���k3tt,,7��y�Kx�쫄؈ɭ�(�E�j�m<{? r�yt�t_m��b�k�� �il���%�1WR��:�ޡ������o��^Z�k堄�<�m���bۧp~)�lr��_��I(@�9�*0���+�͹����Ee�[v��\N��d�~��Gˡ|t� ��a�4�%�#n&*'��p���4�Z����2�%����$J��'>���u����H�%�~�A`t�&8C�%7�d.�˴�b�Z,�+�����ߐҟ8�*/������m�W5X#PE��{�_���}�_[�.��1	7�o�b�_ 1a��lM�m���9��L��A�𧕬m}J��'��v^��*'uӡ���΁\L��w���ݺ��<��=�nP&�(W1v#���ʱ�ќ�7��{�x8/ �D,`-�TNf@�H�0�ܝ�@Y�����G{�M߄ś�B)�P����x��� �ms��g�ΣX_�DM��G*�y����<Z�q�`\F�+���ܱ���0d�2H	<���P'�4K�q�Jڪ�ϩh+ch=����{�Z�M�0	u;Σ^T�I��c�V&�ؐ����n� ~zC{r��k�h��r��vD������T�8�j�^�o���6���Ȇ�}f��1�S�"�6�=m�I�]��WDI0�B�u�B�f2ݙ���S&�o-��h�8�j�
�A"�AD�Ɠ��@s1�409�-�\������2�|��U��Cp5)�N�+��my�L|K�b,[;�M�I`�mѫ��z���d������L��*�?t���Q�$���R(�vqp
7ET/;I2��ڛ�H@o�dy)���&�}ؗ�0�r7��/h���K��h�M{j���������� 0��ý��6�F	K�E��{�����>.���$���?����d�R���x�U���py�N?,[�i!�� o�ѻ��U�����I��J���H�<����@5|
/���#��Ƙ����2�ԅ9����4��ڒ����9�]�������̹���n�a�d��E�"�$����ϭ�'�D�h�uA�ƙC6�y;�!Req��qT�Ga%��;L�L�w�|�X��:���?���|�X�B����V��緘1����xN�1Cn�^���MN�;��`���a�jWx[s�l��i�i��Ë�jˈ�i៘�U�05&V(b�9�,��\�X��Z���D���3Z^L2�z�&1L����$�Mq��d�������Ƭ~�@�r��!�5�!V����_N����+��U&\�����
t�kȕ�
Tt��E>��,v���;�q�v7��	햜2q�}��eg�H��������ZP���Q��E³���{ᄤU��')wN��8�g1g��`�YX�v]&� ɮ��Z��in��W�:�)�)����]>a�p��ystN}T�L�&%�I6Z��}���_�&��h�1,��f��� <V�6Su�z�b�kҧ��*o/T��O���c.�� �k��z�ђ�D���Y��~��W5�����ڵ����	�# �d�FCi�2x;�h':�O����
IKX��Ag5v��I}0]�3�i
0ߤR����=�1]�`p��/��~��c��j\P�ux�2�mh���/��뀽Ddp�`n����B���}������
��6x�+�"���=�g䗔�7+��=A
�<wZ�7[84
y�P�r,C98V����޾r�s.,�Y|���G��.� :�E���i:~7��ܯ'���W�;W���lZ:�s��(�C8�G���\�ky*�vش� �qv�%� �v��xSW�t��_E����"y�Э���5�� f:'�Nl.�����S	XZ����h!4�kbbMԶ*Un��(W�5o_@*@��^�ER�WO޾����� BJj�[~���:�=��A�$��75�9wǋ��eǸ�1Z��F�Mܤ� >�C4 �Եr]I��:o\|���XR!	��4�M.��(��˺ӎx��_���_� �ht��[�M�(G����-�vpk�7�ĉ��ݔs�iJ�X��[�7|�c[aqk�.�Oja��A�CW���l~�I�p��,Sv}�_�J�����UJ����ya�q��e&�t�<���,;^�a�o|<�T�8�#�g��d��/=�>`!#�u;���9v{g�%�`��DO��քd�������<�%Ԏ�[4ͧ�1E��¿B��`]��e¢aA����d#O��}q��MDQr�`|�>ǻ��_%��{j`�(���~��˛ow޻�����h����>Z��4kL,����щ��4�C���#B�A���6,���~Fa��#�9)
��hyBo9��JF�'�r
�R7w�4/]@�%/���ܨ���Q�׳�{�-H�S�9e�9�@q�i{~���
g��2�ږ0m���� �]Jh%z-j�^R��%6z�U���3���U}�ƣn��B9XܗX��J��Lӫ�rS �_h����nS�s	(i�M��A�A:�B����<�qW����/vY��������O&���~�$ �xz�6�
1�}yJ�����ړ4�K �<l��4�y��},�0��,�SZ������_��/Bwj�^"2�~��|L�Ҡ�'�EY�ȧ�E(墇(Z�[�V��'l-8'g�2:�X[��X�[��W*q��KW�Ҝ��轴C�ɔM.�FH��K�.]n�$��uxW��jk��ɝ�������ף���w�(j0��h�j8r�S�3��O�HZ?&�WsE�\^˲3����?ݦ����)�x��Ī1!�7	-�8M.l�0��a�^R~ksY.�G��E��RcE���]�ɹ�.23��̋�G��]o�c�q�r�0+�� ~��>��/-��j���
7����n0���C�ƦC���t���=�0�ŉ������X�[fc=�(�ŵ�{�K�]Y��q$����|9�����=N�:�ca���N���Y�lݞ�ĵ���$������/�8�\�F�F"X��Wާ�%� 1	L�������w���u���[ܴ�:�n �I|��(��T��*�o���1>1B���������vi��
-�h�|P㕽o�u���2�=�p��؍���?`-T��x�qJ��0T��ԉG@2?Dʊ���SCfԿ������y��Ȍm4J�\��� )�Z����^<f��O�xkc�$+�!Lo�o�a�e�'U�����P��ZǗ�p���P2���y���=�[��D{&�%(^����J֠�L(��
6�8>�	[�/�n�rQ� iw4��%�P+8�>_�Ǆ�[{�dk�
ed|�So.����px����d)@>�a�p�@lT7.�����u�������Ȍf����wF��45������y�͆�3�<�W����p��V�yyYQ���H�j�OBר
���_���]��V
�2&�ӻл$l�>����Z�f��nRe�����x���Z���^S�gv����(Q���b�엧�ދo��(�;C�?�<��r�0�O���nmY�K|���i�m�bn�(�L�G�4���^���k#�J������B5�����%oiC�=�uh�Y�-���k�R��R�;{���~��ru�;�s�tD������Z�,5�xT���k?����t>�����`ؼ�v��/f���.a�3J�m�c���\�����Dg��Xm�~"(\9Q1��]���2<E�f����R��������?C>b'd�[�=�淋�k��O��:V����b�W9���&ԓ}J�=Ao��ё�Q�@�G�����A�FN�GE�2H�[.o�į�,��ݕv�,�ܕ/v��Rxb�7_���/�F-�8z�c3N����u�]A_<!0+(�!c!3B8���4 Jy�r�=d,�?St�F(��fi7�Q���`�����K�=��q��+8||��+S���7�Ҿ��z��Q�(AҚV��:��k��^���n�6�|6waN�b�rDB�=�swY�;�PE����YF��.�5�S�;�̡�[��RC�D��p�f��7Q=E���q ({I5����O���<!�r+'^} c˘�e��48����ra�L�Eu4��[���D9u|�b���Fvӥ�^�ʒ�(�̷�i=R�d1G��m�5�N�|��x�z��q�I(��h��?"�
��wƸ1{�24�%�b�8-@�~��CXO�l�r�߯�"}��(�͕b�z��1B|TE\7G�xƮŬAJa>A�nt�}h@���bԔN���ǣ��Y�u�B��8��$�<�T�K?P�q����Lz#��<A@p�A*�r��(�w�:�����q��� 5"�`�eڵ�8��7"��[���3�0È�h�)�-D?�����]$Cװ������>K��\�c�� �x=b|Hu��qP���ƀ�O�2�6�=�������ڤ�9������=ё	)Sr�R5	�g(o�=f��~-x�p;S�f��P����i:����^�ι�'�כ��L�lO&7C����\Qn�+P_l�c��$ruA��|�Ϯ�JY�P�Owh���j�nn���}���{%z�$�S���iǸ�0�������2��*8�����ҾQ���e�	�����,`�^N�n&�jil[�,*�Q�����u�.�x�`�9Ë��҉z��Aad*me~����m
�x�h�8��ܰ|����띓����|��Ar�_����X.�,�0�h_�WB鮕%������n����`~ ���y��f7׏�+��wټ��+��k�>�p����"���7V��S�б�BnzN�{�4���&�峭3����� � 6�X�X7�&ejR�웶opX=���@���Bn�eY�������f��ttj����6s��n�c���o�:3L���_�Q����壘&6�д��Y���g��������v�l�/����c��7��"~(��R�NW;����g��@��
� x���A7�S�/(�Щ�y�xڬ&��Xq�C��Ō�u�)�����e "���X�wѝ��/{�$|�X���Jf��Aįb�����ي�f�ev�"�otM�ͫ{�����G��5�7��Q��u�X��Q��2פqI��f�oi�i-�K���

H���4r��-P(�Z����&���k[M�,��g��4R8X�L&j5��Ѯ,Vj)!����9�މ��Mqm����@��V/��x��9ʜ���Y�C
=���w}�Af�AW�����{�(|B���T5���" 7�E�6D�*��7���;x;+ɠ�C"o�?n��m�7O�+�~Q��уp$o�����+����w��H��Xq�no��A�k�'��l�Ud�C.�?�U�`�]{��B$;�	�G��Uy�q�{�73���x$%�dT"͔���g{�܆�g_��@a�&E�t&Lt����B�����x��7�F���`�,\�p�$�Y�0{�zi��_lSL*�,�y����/�-��\bV�����g�q�1 #�!�b����l:�m���b�Մ"H��2�#��=Y����H��#D@[$|~a�x�4W�[I�/�܇�w�b���Ҫ��f��L�ؔ�D!=C&^I����F"洰w�,�xR��+�L�����h�z;�@���ޑ}��9��w�&���da��j�^����J�h��PҸ�*�?�����`ϯ�w�%!�$��Rϧՙ�m�~v�Y. rl=�b���e$�a��;��ˌ�]��:��[x�����:5>�HU���)��a�Kǳ�Mϴ7��O��,&����+ǵ�)[r��ݑ/��6]��,#wy" ��LC�䥋n�$�M�� q�����nu ����Rl���]G7���ofm���&>�O�i��_5���r�6�L��K�G0�'��#)Z�⤄��ׅ�XbU�R	��w�����j��K%�����/ٻò&�?�	P�L�ӈJ���d��Cl<��eCϫL�KM�[�N�Z�����|7��S�*ojhok��!���|csM�giE�»FEBw�l<�2�h��f���<7��9�̓�O���=6iA]	�.gK#\%���+9u�]�km.��W��xy����v��N,f����O嫧�PwAV1��sQ���s� ��Z��(����Xb�0S"�Ū���!W%#����|&8�Ρ�$U�װ'�b�݃$��Bǰ̪����<d~?ahn�|`(��Z͍$��y>��3MNT\�/5_+���]�p��.�4>�1�iϚ>�ú.e��K�g�s�w�?Ŭ��E��'P�����w� �9e��Y�U(,��]I���ӌ�l������k�>i���F�Hy��[��<��/u�+������

���7ؤT^�¸!�'�M�_�����S׫�>�}���/ �fVtX cg�!��Spw���%���>��[��6��&O�CɫU����_��jS��)��qX������tk�y���M�W-A��@�24(T�{DȮ�Omoy|���?V�$^�!�-j#hrg��\j�[Խ�M?�|�O^���VzUPv\�h}�,��|����I��h/��+M�wF-�?����\_#��)�Ba� �FDNm�0$N���J�O�Cf����9#.#/$��=�}fM�rD�
HaA��w�����))ԁX�517��Rݐ��v�K�٥��\@����OL�?������D��*�ׯ�M�^�~pƞ�����g��꧉R���/�C_���])��=��5��cyM��C�[Y�G�8%K��h^��9�*�4�ؖX�6�V�,��9���� x�[$˅�+J��Y��jOu���g��>Y%ިœhD�Z6�k*f}{��ik{Q�z5�ݤ�!���k�����B��.�1�^"��i\'׳���ޯo��a�W��_U�P\.��<'��p1�f�m΃|��=�P�,W�CL��Y��XN����[�	n�Iգ�Y�t�ǯ`9`���L�8�� ��~A��dm3^�u��#�)��� ���;o� �]�S}Y�������\��wk&V݄�q�Tq�R��S��8e�6H���DPXR �П�7����~�;6a��\�H+L<�����1���S�(�'���]�xA��ӫ��͡*f�����-�K=�7��s����c��n.~^b~ـS�R�j;���i&ȉ4�l��h����2|p���C#0���)�W���nZ�V����B?�w�-�̚����6!t��v'�*`X���"`��m�J���Fp�@�ds�C�a ��-9�0<,�J�i����!��guF�K�����NǚB�K>��g0X�����C�&�k�SX�*H���M�C��s�C�=�Ծ#J�y���=
>X]��� (*���2��T�M�9��-�C/yt� �Q�m�9���aH��>�ZbT��h����Za�b��{c���nf��쌲�Y�#r�O;X�1C5��B��9��M�c�RD�M��S#9"���y���.���EP�����Xx\i�8L�Kz3��o|�͌v(_�%s����^��&F:����ULj�S�?�t)�'�f�`��!��=%K��z������Pb3�9p�mDw~��^Sv&�sR��e��~��������1�]�XH~�2��x�����'`E$��A���\#B�(�w��of���S"���)����l g'�a�w��ʺȊJg���_�V�\5��I��n�❝R�ɛ|�@����ZY�V�DK�/����`p`�o���,�����,�:k�P�&����y�+���S����WĀ�U͉��\�&]����0����aJ�f;��JU�2!���g��0���8m��c��f�U#Q.&bk�J��Xi���(��Z{ {��q��lHz_�g�1�n>�ea���d�"�ɬN�C��,�z^���l ��O�]��o���O*�F����%d�H��wx"��(���YS	R)��s�x�4cˮA��C�`;�W@}�y���13�d����r���t�]��6Ԥ�	�!h6>k�r�x��X�ҿ<q�}��,(�q�5�iIp�h�K>#Nj�JwQ$����5��Ksz�x���A�R���6�P��X%.��0K�}�F)�K���tF�ێ�d�i�������%�N��>�K�<�E~m��qc{�A�QrmJs�oRDB���Bu����T��(�˻�4�����@�M
5:��͋8Ibƈ����� �{�l��I;
wQ�~�=쾅'�_^��䚼�P؆�Ig'�l1|��;DW<c@Cj��jlOk��\�=�T{l��ߨ�L䣈Wl�[~���Rlr�#�s��9z����+�c�QE�G�u��t���Ig�?������>����l��m�f5|�,0�5�2�	i��izP]���eS��C��O���	E�/ ͞���Ix��&)(��5D-�N�y땶��Y��U�����0R�Sқ�FOj�Nl\��RJ�ف��?Iq��{I~%q�Xh�����+�ĕ>�iS]�(^������<{��d�cG�{X�g�L	���G�"�H��u�%N?ըtl��ǵO�t����/U��^�����Zh5eѼ>](+ r�ȴ$�}0x�1�&Pm#�q��8U.Z��e?��m�lc�s5ri�n�%�՚7"*���PϿ[ĸ
�Rm���V9m��r��'�2��s"�ĭ�"���R�M�?�>9�>�!�������:�IP�/�O/�xcS���!$.Le�ߩ���[N�Oix�@��ilt`�῎�;��V�^�HM��,���]���<��r����f';�f(r��=��D`O�j�m�"��w|�ңu;�WZ("3� �>oW���l�$Kw/.d�B	?����SI~�-��L�{rC�9ޱ̃z�{S�^���Ah@�ZN��{��+E��t��[i���\�N�^�*�:�\�;	T`�ѦmN������e�S���\t�kE�d�Sua�!<Q�O费व���W;D��jsR�8�L�Q8�<��%S0t5���$�������z8B�1�l�0��K�9")o�w�&�NL�#����]0_�D��!]E߃��k^�l������'G-�;��K��'E���V/2/q!i.����ȤrJw:7E�9[bw�m!�.t+��9��,`�J�/G���G���� x0\���Mz�.�D	���R=�-m��?H�8M�n�A A���I�6\� S+O[1Apn=�į���C.��S,�9g醞[������n�< B�z��YH�x�-��>�߱�z���	��֮tmX��xrm4eA�e���J�JY@Il�u��m�������V��7�r_��(8)ϊ�%�A�p`
�|�2�T�E�0�Wh [rAH)�f�~���~��e��:@�d�OԊ�F�w�%�N�L�(۫�A�U#m=��n�S4`�����lRõo�SWE�pVs�@�q�Lm����t�l20�����}��t��U&3	*�wp�k.���Ağf��+4�mM:�,Q����]@���꒷u�R��~�QJ*�K{�@��-��v�/�����r�������%��--Y{�ħ0-+���0쿸��-~0n���g��K4L�C�����×���������f� 	���� ݣ>��;�����L8��+]M������pPE�;�?$�$|��ݬ�)~s�$��&I:s��y+�<�^�s<�V�9�[!�l��"�
�^Ր�4�&�4f�o���q�,h-����񸌈f�˼���gh�J1����H;r��p@]���Bխ} :�"�Uu˗'s{���AҖ�V���B��P��I ��z��M�V۽����!��	���qU(� � �rq7�s0S�ܽi41V��>^F'k!�U�α��I��E�,�rl�ԅD�"1.�d�����姫���?oM�~2�� ��3�r��Ti!ST{���&���l�Ki�@R_���u���AK8�4�2_u^�wwar�p��f�0�H����F�
�%\#��_u�/����)�5Gʬ7T�P��
�Ώ].��6>�N"���#t��%�2���2*Y ��3���i�6�@�:8>��"�#f�3s�ûV�A�*����u��|��5��t$;�SG@�	@�{� 6)��`��js�3�5��7�`h���?&b�=�3��#��J��~�
=V�`�!�*B!s�Y���JC�R�A��=O;t�rm���1�ݸ�׃��E�$ӥ}� ~�QLψi�����*��8����R����ۙ2ݶ���,�ַ�fA��n0[TmN�3�������Č������p�P�^;n@-���Kc)X'�ٯ�5�E�e�n��T�R1n0l�ՠ0�+�Ca�����@�2X�]��+ۑ�R�4z����ل���tz)_Л��&�Z)�6�O�В����_bƯ��������"��Ue>�
8�ǌ�\��0]|#y=g���P2ra ��)?+�}�{��<��=��LJo�9q�_�[�F����4u_杽Y8/��Cב	<Q� ����:jߞ�~u}���㨍a�V_�S�>nK�[E����ǡ��������Ʉ���6c��ߩ!y%�S��d���_IV�Q�9>�+N2[䟅�>< 11*��O.>tqFx����zBP�cCW��w��SX$/H�lt����̴����kGe]sQ~���U����1�2M��j��\�����]߿N#�֍��ֶjr�ހ�,��Z�M.uX�bL�a�;�b��ɭ<�����X.m_Q�*���"x��L�:�g;'�
D��P·���h�4H�:5v �����{�\�v����U	�H��6�"p]T�|CJ���{�2�(�f��I[Կ�/��BժQ��u���fC�4�"*������ԡ)��H'�fe2�������v���Q��
ʝj_o��D$�p=rdj$��;��2�3|5y�X��r�9��!�=���u�gj�Pټ؍TW�h^�,=o���3��iG�:;��T�vc��E�BO>t5��=���u#���[߶�'Y��Z@��l+�:�Z�Іs<_,�Z�Uk��ﭵW�T\�2]#��&���tr��o��6�W�R����v��X˘�n���2U�#����v6 U�~�M)�2����S_F���B�s#�~�2��|�K�i�f��bS�뀤R?��WO��Oyi+��Z*�?��{͟r�b^x�����[}�#�=����I �J�dq�bT/,�-������P�9����+? v�!8F*�2s�M��Ś@�\H;�3W�_���������5�^���'�]���c'�/��b�p�p����	�U�O'�1���b�$�8�[}x���6�AV!�d���li��~g��L5�r�w��C�B�"�|mG�	ӫ���sЅ�ɋ��w�*�.󥯳�,:A(���w����B+U`
��T�5o��KrʄUj�`��]�~uG��Ӓ�#AI�@^��ˍ��}a��[���m-���~#�x?#�WX���[���NN2�LjwT_n����;m�[�cp��րB�M�/��F��0���WqB9�W�HA��틐�[�!�)H�m�X_N�ו 5%,��}^s���<f�?�� Q �������ٯ�,�� �mE���T~9�^�S������6���@=��sh��?ճ��-��<�)�̫h\u�9��u����W�uLp��. K��GP<,|,L,۾�7Ps
_k|.�)H�NL���^6���O79�D��!? ���п��H��7]f7��.հ�P�;;�ӈ[����E;6<������'6���P4E�FY����ltV�f�"^/E��*P��:�������^B�{h�ex��Q�7��t���j�C�.r����Y33L�O,6P�%h��Wz�#�.�!�lM3őjS�s�����L�Z$X�]c$�_�ja���1�?��,��%��q}Pb3H�K�%���뷩41fB�[��ŪSё�+�G���(���P(��X��6�I�:r0Rd-{��5�±p��&�>Ȱ�$EL����@a��ۂ؋]LL�o��{�Z�w��l��������!�R�{
n�{�jP���ݶ��[>X
E�,��֩mu�؏�	����	u�9�ф�Дר	�9�fRo�>���6�?�x���K5.^ٞ �<�H3U.��}ԁ���[Ү�1�"%#k�m��Ut��VЉ�{��^��i<*���);�.WՊ��~��l�XT�3A����y�(`k��le��i�z!~X�Q���y�8JcN
[��QNO�L�Tմ���+�g��b_H8�(kء��?��_}`f��+q�� #q��-E$��є���U��Stti�$��2�ĭ�(�C-���^���˵�A}`�/��� �a��Y�٠c;PM�ud�, g"��P���}�)�<�U����z������.���]�"���s��A���\���b�3*
(���_
�z��$5�6/�Ty9����tH1������I�'��x�[~i�lg�W�M<-Cfq��Y�Cn0�
'{ ��"�i�ZB�u���5O�6�J�0z�.=�<Z|݊S�nH�u䃥��b��$�j6��r9���&�qaR�'���VW��#�H�v����DձG�s%���.�@Z��b_��#2��	rbm���c���������6h��\Ly	)+ ����Ss+�>���K�$��	�-BV; S��J1`���E}��˃���_v�T%��W��0�d0@KNQ�1>T�ACG�n�U�F<tu��vR�qHb�\d�4��Z���r�ΰO�x�nYp�n�e��X* 8�L�EB7y��CV ���`�A�*�XT������ͫcg��^���ئl�-y�?�H�]��D���e�\tcn�*���ǰĀ.&�����f�m�+���.-����B��Q8��O�W�*ȏGЏqw=�.��!��Yܤ�[��P�Z��q�뤢R �"�uy��B�o&��°�
FY��ܷT������&w�����Hl��$�*�����$aqB��n
0
��Ô����iZ���	<�h�,��a�t� ��&�u�$Go9�ﬣ��^�փ;�ǉz�ή+�[	۞��R�Ӹ�þ����3���2�w�}��n�u�J:����pÐ�c��u����x"EK;&	y�f�Ui��}���o�� Qw�]��%��)�8uKyqe%���E��)ۖ�'�����F�1�h/���ݞff���F_��ѻ�Ah�������Ē����Ƕ\հ�^Ri��&�]~�.��42����4ـݶ �A~N��<��y]���O�.{�������("��/���ouF�AV"\h�۷ �z���#��2?Y��X+=����ح�Ia������_�T���Wb6�-�==��c��\���K.����6Uz���F��"Fg�:S�O��G�W�}���Z��荁�m���!	��v4��&�v�n�$�x,����̠�]2��K���e*��2!�D�Nu���u�E���S�͔)�@�ˑ4�L�-0����N�ܠ��tSX��[b�Tj,�U7��U}Kl(0��d;���l������I���'ѰQF��J4Q!�����5����j�[X��0���1�^�}A�=&?����a�֐	S���T�P�΅�E/.����m���,�q��fX"�!����HYe,р���w]���A��5�9�qA�-?K��B������!6����O&���wC<N��\���N�v�&�L�ʟI6�@C�a�-��!�b��d�:���h�ݗ�%w����e;j���rB����#O>PRO.cC�gi����H��s���d��(���U��B�B���e*O܈SO��|0� � ),\g�H	#��S�NMԗ�r�B2��)#�$�p6�3������{�91�_>Lp����ϔ��jI�E�@�S�r��
��c7�:��b�-�o�,��w~�"�̀L���^P�h��â�c$����� � �f���n�P�΃B�@���,�v�ݏ��-��N@v�=K�&iy;Q��`I-Y��>̎�����Å��
�}�$<<��5}�,���*9�b�#�������Č���Cp{	z��?\ehz�z�!��s�^f�I�����*�7����S�W�pS8�f�-
�e���Z�F0�C�7��K�K�bhv�k�V	j�E3������w<�W
y�1�9ϛP䷽GT��:=ma�3��K�|�]`�Ǿ�"��n���&�ӡ���>��^�sys���ǲ��R@N�<3���gg��&��G=J����桢��Ǌ׼��	qߧ"1mS>���t��Kt:/�~��aN���<�v�p��`�Ld^��w`:�����y!'�����Z[s�9"<�e��cZ��Gs�4y��HM1��F�� �<T�ؓi����(�<��c;OR�̤lb�(d�
�EY��^��,. g�ڳY'����w�W�ׂ�?w�8̓1�ۿ?B�J��n�45��"3e�:��&�P�ؿw-��W\���k!�W��V���m����N��[�����v��ds/���Y�V!.�˦��V���܁�}�иfW��3�U�+�^GE����>�B��-�³Ӕ��rJ=,n�+}�V7#<��5�f�#v8 ��vX��e&��J����T�d]>X�(�gbm�i^�V<�Ӫ�{���fV��*�1�vԋ�P}k��+�����`?RhO��&$~�}�|��b	%u�^~�#G�ΒLf�3~�R<|�u��.���R)��Z�ij�	�*D�Y\a������~ё�o����n�?�Ժ��@�T����]�6	H~5y����n�t&'�M[�f2e����٭��շ��J�o���(��?K�eQ��>�*�R���@a�iw��A�)��J��G�g�S0	���5|����筫�4�#�_���Mb�=*!���[^^��I�,�Oee�%���*�zZ7W��$j�M3~��W�e7�QU[zt����HK=E�_�b�2��Be!X.i��xU�>\��ʹ��|���>!�&��8�4��0�)�O�B�	]
�l�w$�|S�h�Em��:���������l��.�U r��V�h�|6�S�TG��LƄq������$��W=]�i�z(ĤTV{_~'a�m3�r�?A��WVE��aOݤ�q?n}�F�h�炠F&=PL��lXqF�ؼKp�7�P�{V j	�aV�:�~)��y�C���7�����/�%V�a4XK0J��X�aOk�G������j���Æ�n�j؜�{�����j響� ��4���7�r��k���Л�x��頁L^9#E��_���Lo�P��u�.�^gi�̖�s��cַ��#Y���lV$���b붫�{*����GL0Y�
}t�O��"��&V=��8
��]=-�\:�F9�.�P��(�i֛��{o����SK�M�w1;SڨJ�J"e��~�>u��=����(�=d�S-��i�T��I��l#�L,�@��e��X�[�j!`4�W�$O���RRT±׾ �uf�*%Ug��V�$Rx��k�a�&��O�$���[�O��-�z�L�N9{�v<��`�ﶛ�_�(�	��t���ա��f�+烥����#mކ��|{�-�DF��&�N1NC�==��]Re�H/7���'�擈gx�!*�&7U����@	����q����f�91���C�&͇=� e����Ū�.k_ɾ�PW_͏���1*�sP,��~�Ό�څ?X�������:�Y����}��,<��"��9�q(��n�dW�Hh���A"#����w3e5��!ߋ�����d��+����ut����
*�K��>��,���)��<O��z��VSWU�$��W�������w7[�5u.��̐w!x�h��� 6�Os�q�^����J/�=�6����5���g��$stâ�����s��L��-9u��Y��*�S�n�|P=0$4>����Xsf�W�k+��
T�@���\,&J�� ���$�\0���.��Ū���60?$�!(̯���[[)�:|��K�8\9�����"BH��Gv�?�K�]u"3D,��7���Ƹ�ɭ�2ˉ�}rz;XU�[��G�8]0����ГE}T��v���+c�3��Ԋ����<�o�������m���?MV �p�(���cL�?�]*4-��_�x@	�v�HVݕ<?��g [�ǊǇc1
�H���F4=�D�#Z�Uѹ�'�Pk�P�� W��8zx[��-�Q~�M���Sח}�M"q0=�ƈ�)��Ck2%��Y�� ������T�yF5��^�>wt�*Q�����<Ga���AEDrM�=�q]��yci���0�aZ�=��rc�v_ӻ�\�~],M
%Xv�B��~{XU(7�=t\��v�T������)�L�_���G3络�O|����:Q���O�͔��Q-)���\�W-I�U�+B[��?�[Ք(� 9�5K,�k��1#�3�Ҥ<�"�Bh�����I���N��Wy]�f�� ��k��a���{�+���Bt�(Wx�#ʙw�>=�c�s������^��ad�:$��Z휫�m�l��'L�H2�7�n,��M�N	h��{��I�M�_ј�e�7�Lc�L��觨ݛz`��A\gNv�%^f/�>G�x���&=�d��~�vq͝|,��1�J9:O��b,}Ζ��x-�)!�XD�-�Հ�B���WM��@�z�35s��x$�#����۾ C*��Y��˪6����*�O�f����c��ſ�0�z0���Z��:aa�>*Sq?5����`��y=��ɩt<&iUf�MA,H .ʨ���4${N{��2Z�bJH��`�j^\�Ӂ!Ӥ�Ɂ�/��*z��^:R~E2Y�R�ھS~�EX��bz�?�'@��푠NVx�7\mIx2����p�{������6�(��4r��+�oV�s�=$��V� ���W)���%���'�sg�YuEc؛��`�;�e��yD��1fx�>5�6}�"3�L�6��#K���w�T9���l�?x�}.�
t�Va/i|�t�Uwo?�����P�r,�O�`���b4Sg]#����l��n A�l2���O�/����&�yڤ�6�3VȞ� 3%%&=�_�3�z���
��'�=/<77��U�x�� �Hq�b����{#$�lAk�k�E1��ٯ��ؿ$�n)��S0"��U���A�á�T�X7p*o���є�%w����h,��	��/���!��WP��K��q�0��=)�褏#�x�%d�`�����K�����-�N_L\�*?� �.%7�?ќe��ܟ��湃oX���w˦���k��Z����*�gژ4ޟ�g
�@��������荫WP�z���~�����R������Nݎ�cs�ׇ4�5�0�ƥ��f�)�"©}�����V_���Ș�DCB"�����M��|Z���~p$NƖB�^�˟~�-�֙����ށ����!����s8�J���mcqe�P���& \1-��<fj炟-d��Թ�WE��N,_b������H��7�J�j߄y���I�Qew��1�-�8�*;���zZA�tE��Rf��?"�h��tY�q��F���(j��wɼ z`� "uH���ǿC���/C��/OX����Zg��(��m�ђVD��R R�(�1�&��p8IP�	<�J9-�{��}�=z٪�u��%G���pj����ڰA%3``�)�|��f���%B��̟���8�j�L��M������ J�o&���5��X�S)�0g:郰�� ��� ��ܓ�$:�߽Z��y2�@ca!����e���l�ڌ��/?�ZdG�[�d8�bSUt/�Y�H�A�1
��W�X��4^Lۣ�Y�6@%Rpv ��q�m
�!De���[\G�C���U�C����(>:�!�DB?��Mr����	]�M��8����> ������W���:�Dĭ��YoY&�'g��'8�J��� �$�����S�&����@�5K������:�#���<~�K�U��}�$�W$k�-wׄ������|˝ﰺ��j��L\I�
n��T ��p��� ��S�3�>�W�G^#=�0��.��/h�� N��\w��	��[z�[�X�,��ͫ<ğ�&�<�M��We�5���Ad	�U��b�]�)�ߡ���_|[l`��Jpg�,���BqJ�D,�XEʤ�>�T�'���,�Gr�jlr�S��]vX]b�a�)��]�R��k��S�_oi��lV� ����Ӣ��;!�E����,X��f��Q
���-�9㷬-l�v	�U�ſ�;T.�
��/�\�ŹgU+Q]����]QK�ȏ]#ox&��8��Y��$#�SO�uS؁�N~�B�/�H	�1(i�I�Nl��<bcpTv>�P�<�b8�	lg�+�ź���f�e�7��;���)PU(��6��]�|>����'a�
C6S�=�`�$5YU�X��c0�b��ޑ����)���@|��ܶ�XFON��~��$��i�O9�Ѿ���X\aע��,[�6r��	D������V�B
�L_g|P0���Qt����*�-z����|1)���i�׸|z�_wA}�q�����~�b�Q�M�oʞt�Fˬ�_.��h���oZo!���DZ�(}�S�[мx�]��~�JB��3
���1Y���#}�,�l�N��U#�Z�ޙM�(�C�bC5�ִg~�i�	�rARw�ِ&.@sU2���̕8P&%Cu��5�N��L�:����4]��Gm'�50������'�Rj}TJ�� ���2*{���QD����c�V9	���&���kX�&�iF�&�z>7�B}��0�ߌ�e:�J�X8��U���\ʗd�-�*���ٹ\}��2R.狒JH�]Ssln�/Ƿ���r��"�Ɂ���y��5S ��m����*���?ƔS\�dE��Ɯu�ih��W_�%խ�yM��"0�T�<i��0�g����y���W;S�Z�Ё�g�|G����C�Y4���c�U7	������+��9r��I���NZoͯ�rS8��g=�<�����K�8=q �Z4��i�V����*��nG�	��^�~�S�.��׾��:k��}�
x=����E�`�V�N�PZvMi��{�+y��;��Jie�]2�O8�+���3#42�?p+��lח�:Oe�2𹏖�[�j\�����������=F8zp$��>G���T�Hb��ӳ��;��@d
+Q!��_��x!@h9JP�!U��kK�����ɭ#�w˴Z����.x|�-��W�P��z��K?�k��ܻ<������6��!"��ڬ!mA8�3��94�,��&�n����My�g���؍�C�3Jo�f���iKz@�	F�!�Y�����z@�-���4�4az�?�8��2��*�R�R��u�V�$H,�޷�����3It�Pz����^s^1��ui���<�����6��n��x=�e��)��[R��SV#�ryJREU�9v��a�����7Ƭ�u�bw3������I�۾=E(U���I�luk���U���*��h�e:G�n�q���$�Xo2�L�������9�'���@fШ=3+\�Mme�M��E�[(��β����G��b)�3t1Ӭ6���+���Z���H���Tqn	�$�(����hh!5sI�����2h3�wQ�5a΍wb���~�u�X!̗Y����^<�@mO�箠��@I�H��9�\�G��Vc�j��	Y�Q�.=y��
��_g:���{y��ge�'![�_�<B���z��<m��^�{A���tF�;�T~3c/cHY��1~���݅8���g���wB�1,�tͥB�\yȈ⋑�D��䘩p)6��� ���{��nw ��D�Q�l�w���۔���e�}��e"-uY�M�!f��%C���x�e�y�������Q��ӣ�u��Y���i&��g��:ԡ>���\�����
�~Aa��~i�Mjg�`'/b�N>}sH��T�[�J=��_�Y� �0�}��7�F%��gg�;Y7��P��{$&z@	��YS�����پ��I[XFnC'b��d�6�vB�{褆X�By4�m-a�NN���^�w���`�U�ws��KTq�
e��=tMٶ<�A�m��DVu�zU�HFG��G%f�I˺& \9�[��x��������J/-:L��o>�6�+\!r+@��k�C^�<鑹�Ig*]�o��At�y@�f�z�0O�cA֢$�q@���u�;aX� 
{U+�\[�몰�WKx����lm�����ԗ����f�FC�W?u�&��ۉ�lW�c�룙R=�ߴ���:-����-Sl���������v�T���B4j���;!�:r��E���\#��ʔ�PZ��q���L�V�Ȗ|�?Q�B%3F�GpE��c�u����&��?)�e��/���vV��Łv�sҸ0)hH	?Z����qol_�(���l�� ^h%���ܰN��^���=�V��H=����2�W\fs8�l-�*�.a�Z����P�;�Kx�}_G��CV@2s(s4O9l�r�oӨ�M>K���)�r�bյ��-���[��\Y���x�y��:Zu�aF3�J[.!��279�}�8o��Q�bֳ�ơD��IEqLs�y\L�c����l�9~�ܑg�	,��h�yӥn� ų����$X����Oz�Q�rc��4t�+�%"��|Ց.��Ͳ.����\�@���d�"WT��-~�-Pf76�O��k[�ǳ?�zL���ٞ���?�{��)ײFҘ`��a�H%�c�C.�����Q�\A�p���t�C�h u\�|�vbHҒN�a�.z=*��g�F�M��(ɣ�\� �9  (�������� Qy��������9�z���{��w8e�幕dI���q%�B ��h�l?]���L�&gI܇P�ݼ��J^q�!@��6���i�_����
5�N�&�4���Um�&�#q��14˸�G�QQ�P�
+�- C)�P�&�;�ii�^S�b>����\S��t�`Je3�ؔ%�e��rsd�`�Lj��$F��+�8p,����z�ws�v�OZE�1�	c�-/E��+ .XcO)�/�$�̍��QW���ɶ�_�l�	nkOa�OAR���;U/�Ӛ\��R24f�J���P�Ug�������ɥF�	��amsR..̑��w�7_�iP"��F���U��q��3�?l�_[x=M�^�k�!Z�7ߤ��&`��r�Z;j	{�����B�Xw3�F
hC��_H3 z����}���#�\���	ѱC���ׯ9� �߭z�����f�8�a57�R���@r;���>�-R�𜗞;ƣ�����?/�f�$�-�����{~u���y��[n�r�X�e��'�����ZQT�=�r�x�q+�櫗�deTBƯ(�����\]>ury��`�񹔮!�{L��7^�_��3�����9�eڱ	�];4�lo�h1�������^��}���Ib]UT�T��K����zw����h:���(�?	�/���P0�Zp�cEv+=Opl߂��9JV����|��mATɩc��f�V�cI6��U,��>Y�>|�`!���QO�����qƼ�2	� :e�4:m�� ���l#�C����	�`��r����7��!�\��$�)Ǽ�"o&'���&l��t ��Z�mh�Z�Z 4�����.g���)2y�F%�4�Cɇ���!m!w���$=����d���5h���e\�����wi�)Q�l:��G~�릛0�
_�t�2f(N�Lf���m��	,wֽR��+��ۿbƁ�c��`)S|�+:E��Y4=n�����+����T����+3�Ib�Φ���ڃ0�+�o�������?�E�(e��G�B��:灣[XY�<`I+�
�[]S�ŵ~��I9G�$V4;z��P�D�
>IE.
"�|��
�#�c%6�rM�)��,�{)�FB�� �Ķ�����%�7.9.��O�ej���|����a�?�U�G���.���r��ɐ�����8�*�)E�J�����m}�Ï��߁���n	�c\�>��]���[HG�y����3�ǯY��_Dc/�Eց.��Ҧ�j�h��U�:2�#7�$�!`��)r�F�9��W<tv2C }A����8���mי�g)n�lm�������$>�b\�S�T���{������vD.�t��R�G�Pp��E�e7��g�c)�5to$�p����ǮI��3E�-$�m����^U�l���P;i������E��}�Y����ٞ�^� [A抸�f.��j��+J����aֱ,�Lg�7Y��|�����%����7rb��zz���t~=g�뾿�M�E2��qhQ�ڝ�?96k�<$N\s#?�,�D��z,���w1S��ZN��w�и�;��yed��(��@��~��c�]G�c��]���Ȯ8|,�؋�:���;��,�@\�Jf$a�F ��������>�z�Q�����s�S�_�%y�N�<���Xo�
ȇϓ�����|�%6�n����|���V۷�����.jj����
�	������'B!����C��[�UP�?���a���8���-���m������8S����U��@�Dja�I���V�����-�)'��%?�E�զx]l��Lۋ(Sm���� �A"u��O
$��*1�Ȧ{w�"j����l�hU��hni޽lw)!j�.��(��N��3o�y����o�+:�F�"�8s��C��$��6�����fs�h����!��|yBQ�;�&�0�U��;��Q(딫���b�J
Kuf[,b�ڞ π Hۿ�X����j��7RSDs��l�HmMpf����	+�iB�2x����Qn��][�`�,٦���\�@�R Eo��xPQ�`�����̣E*n�J;�@� &���G,��y�{�:�*�}�k!��ﭜ��>��ƓU�f����5MU;7�R�WJ��E�Zq0w@���L�H�p�4�A�硴tW\PHH
��큊O��ZM��Zo�����xN�	�'����g���-������G[�& �L��Yg�q�
6�R��Kpcfg��9�&�L1�<m�h���ax���_�_�׃dȷ3i�8G�B��<1ώ�1��r��C%*������I��W
3*�� 4XD�/f�Y7o�I"=��BbaD����"Ռ*ml:���n���ԋ}�؏�;�[(lYW�$M�)�y,���#!�3�ϵk�c����4��4��d�I�ޘWM��ۡ4���H>x}֜�_K}Ѩ&J��&z0Jڇw�r�OyֱԵ5`�&QxIe ��8�(0��0����,~p��W���vv�Tt�JK�ף^`��L�r-��=jx�N���Tj���d�r��<]�/j9l�E����1�qE&f��T�GoM�Ч��F����X���݅F�^���J뙎��V c�po�+Da���l��Qw#xD�j��;Ƿ�zJ��5�>�7�)`+���%�@����$�����L&���[�@��-��f�G8}�1�����ti����5݈ ��f�G�����ɨQN��V�b��YYM��W͟�d�_��`�%��g��󲷄Q��U��u�ı�/8�`�y�Z2�S������;sYم�hL ⍨��m�A��\�M�_ǐS���@-�d/#���+�u�071 gMR�������2�b�m!i����?�V��k�����9�pG4^�,�)z��Ey|=�AT5��-=�؅0��b�_Q��خ@ȫ⽒̱XL�hݑ�x�_~	���l��:E@��`��7��� ���e�';����C��`Ԫ���\�w�̟͌ |�P�`�T}���:A�`�ޣ���|����p��hm��?��(�M�A�J����('�� �HxR�r���oi�� �����N�t�ԁ��i������ߟ���i;�n�c�/P|���/�&5Ӣ��(�����(%���V�c�
? 1�n>�k�@�cS��o�1<��z��㐩˕��	��h}h�^	�+�F�����~�
��3íORmV�=V+b��#�Rβ��f�6~ōI-|��i�G×�PА��,�i�i���{E����?�r8�����x�`l|�xo�$7֭�Nx�e���~�W9 ,�gU�#[݆�9���d�;*�sT-���U&�L,в*<�)�bk���Z��h�s�6  ���3A'�z��H�V;9�#�.ym�����H�QN)xx<��բV��֝�޿��������m��/�a6�9%x�\�,I�����-�r@E��ƀ8h9u�CX���;^�O�O���{-}��3Ș�گ��w�G�X�h=/��d�f���৚W7R�#������L������ �j��,�@���o9Z���$}���utډ��X�D�tA�p������M3V��D��#�'�Z�֜�s�{1sX6B�_��ϓE5�&�({(����)��C����{q>FoV�M`\P9���	|�A�'��������U���Q�(v�nLį��9�������r��َ��V���b��M�s���]	A��nu�:��e<�t:a���j;�f�81K���j�x����b8�|E�y+s����-m��İ�c֧��Sy"@�f�����3R���_��]Fj:��j��]Ϯ��>�Ш�$ƌ�*��Ũ�r�o�.w��5,o��h�#"X3O	w�D[�\�Bjk�QZ���@"�6���hM��@O�'S����{I�2h��� �������_�܆r����.$2���� �:㊻��6dNC�g
�����`�j�����t���s�v�j�{P���3)��(�6'�Py�Z)U����Pc���P���K�tZ�d���ߥZ"
~�
g��[_e���9�{��_#@�����0X��	��
-�J���#_�6��ܾ�qn� ������e�X�(�ˢ��ܖ0xB�Wݨ��El���S�e|Nyō������n�Jt��v/���5��nF�3�B�9f�d�ݘ��_���K�^BeR���$����D#Jz�hQP�$[��+�|����0�O�1)��삫Y�����T�8��O3ܺ�Y�	��N0B��DԼ��<��q��c��m���	�Z;�J����ҟ��W��}��0����Yf�3�z��!�sI�q.�m?��G �_�g,��E�[�U��gu��n���#q���� ���?t� m�_�,ILLW���.�]P�4�eV<�
]�<Z���D����Бb��=��?�]Q���`f������{�8��ERC���4t� 0ܐ����
���nF����\FA��t�V��.�8�=��#T1���*M��@�(�\ 	�%)1�:���'?��<�[���$!�@�'Ӓ�4nd!��Ѡܖ�Yc}*��s�6n�j;Ə;�����5���!��K[�,�4�|G�������r�1��%�Ovx�������v�I��p|�:��+�8�*F��lk�/�e��ˑnA�%}J���Xyퟸ���g!~�?r*�"�w70R��[9�Џ*�W��dM�u�%��Ajð���{���ygf��1�1B:�������	*A�T��BrңGЯpH�HUK-����GB�s�>Y�j���&_^�3���QY	���r/�Tg������}O3㡓�K�p�i�ı~��	RU.��V��а�9a&�P�Ș���]lEu@��T���9	 �6�'�_7t�)=SAL�b�lT��R�`G.����u�>�H�,b�?.�V+� �t@�K����	��O��H���=��ZOJ���#��z�*��&`Y7�?�v�X�i���q�a��G����&E��!"�ϭz@{�m�S�Lp)=��z�Ğ���#��^GW��=��K%/����<��|�J��N�1�:��`����%�=�7@���!,:�>=��3ȫ���j��66��� >g���F~d�Ĝ�b�en����RjE���R�����E"%-1zDf^�cl�[%~�є$�4p�9[\��VM�:*
@?&��G���2{�����P��6��r7��q U �E��o|"d&����Na	�q�K#��p�~�OE���=/(p��"��t�&5�����@�Vx�ffg�ZU`�W�\7�M{ؙM\��퐯�k ����>�bh5N�|�X��:���%��9��&Ф�߆���eYkq�,
�^��Fv�ec�0��(�a��z���\�k"wj��������m��i��H��%�tc�j�,�7+	�������������SzRDv�3;$ ��q9�U[`��k}A�!�un�~�
����z��:��X��Kw~FK�,WC%Ox�f��^K��Oi1��3gP��%�
 g}�y�/q���G+��>�nwL���X���	rbB�휲_��oWBX����eT'��:X���H����z�����ܪqQ�^BGKL�!>��C�B�(�ۗ۠�����%b��>,�q����Z�x��}O1�s]�-�.x��<�O!��F�gN��}C�K�g�#)�I���ߍ�Uhg���:ҽؿ����K��(�cb0���C�da"8�^�h���
l29�OYc��_%��/�VLݭK�0���F��D����1�\�m�e��f��T��"��]e���9qޚq�����F>х9S�
�)FG����.��?��L\�ש�!]��(�48��eR�Fy�����S�"��@K�d�Yj:���X1�_��k�������=�.��W������h�p�yM#�>1����W�+	�5c�Lh�B{g��S�Ԏ����M�¢|a�� !>n\r��ML.ҒƅTf���8���Ei?	�L����$G����e�ا���-ۖi�%䡣R�k;:��/��P��.�P)94*�b;��}�;���_�|�%��]�}�X��"(���/Xu��T��)̽�"��	�Ό�?{��X#�Rds�ѷ��`�6���62��CL�O��$PB�U׎����T]��B$e�o������G�C��0;	3���6��pe�jپ����.]bׇ�+nj��0	����nM+nP�< /����5���B���t��4ww9K�X�Tje�p��z���W��l��x�B�1~� -�V8�Zc�2���A'��,�����Em�^$��n�D�B�K�4�ac�F��6c�w���Z;�R"э��uŸS���̠�t+Ѳ��h6��+�Ƌ
e�Ŧ�ݾ��|�xY g�0�+]T��6B�5�/�͑U�JA��i-P�u��:���2@�#{*�&%/��yE+"r�$p�Ï�^�7�T�&S�u
�=��b����=ìH�C\�M������]�|r�� ip$����pϲS����$��B:����\زz��� �ש�=�?�V#ԋ��\�/���o��&F��x�ƶ���e�c+&y�h1���*�.�kӁ*�Yx��A���Q(�!�hf��_q�|�į9��R���yˑ��[u3v�-O�G��{챪���PE��:n���=�����4�o�Ѿ�;�:!	F������ũ{�ݳ9x��<E�@�h�w���2<cYٯ����
�x��Ie��G=��I�ݞ��=l�"�mR�<ۊ����s����y�/7�Ġ���O��T��M�pF�$޿g���w!��]��4���o�'�[3�+�n�J ��'j��<�c)�ǪR��~:��k/�a�)[����^6�iN�PM`�ߍ���5h�_��^�f��`�M������ּ�
Ѳbp�,_�lCnD�^D���qw4L1�a�'`�)N�:[i���>U�=2�I�B��vKqm��,*f��K�����=sf0Ґ�#8��Fd/BG��y�K	Y���Q�x�b���H�cr_���;��X�۽2�O����r�����Q�[�s���EW�a`�r�Z#�f.�\:�|��D*BR<�4J��8S6@oL����-¾n!�:�["�[+\@��F�>�vǧE%��s��_�L���s`5����,�|YR�TX�q,��v�ǽ{ݶ,q%|�_��y]ҢV���M�Y��.�L�\�fv��){�m���fhTJ��9!�� ��qD����b֠��"R�����!PN�贯CO�f�c�{���P1��&aS��/h})�+{o����ojY,�3��b�����eʡ��i���=�M��7fa�dqh�mo�h�它A�p�Y1����<X�>��'庒�e$�{�x���l��Z ��C��Lᓲ�t��H��`A�sY���T���ڿ,	mB�wE>�I)�DA1���9�ʒf��ud[���aS#1���#?D��z�-�'�N���./x��'�!�J��-l��@mj30Ω�_�ek��cZi��p�B�G7d��6\��+FY���[01��ľ#,��6�x+��g!�e�m�m?�>��v���{��ܺ�Ԃyn�SKV��c�ɨ'1E�$Z�aS7DS\�F�Y	�s���ZA�CU9� ���#�i)KEU\j^��_���1�7�7�=P�"�@�BVx4(�f~؎���R��0�����c2o}~�[<k)�q}\�[^��\���ŨM�t��;������# k�B��k���������� ��;W53�|l<��@�si�Q{r>b�^��p�V�Đ�Wrc�
+���t��+Z5�F���[���;��_����]�ܡ�Јam��RI�V
B����NT!�E��sX���Aۦ�(�e�G��" �k�T��C���X�9�E����b[P6Z|�.�TV���>]-s"K��
1:)��+̶:΃B�]�.��>Iϔį��@�l�:-�-����5X������w#s���wV��`���Q�5���~���6�HL
���a�H���F�̉�
��c)ڃ��\0��N�fjy��jj��v�0_W�v#���Q�sr�]�f�A>�>b;W�WWΠ��=}_��a�^�u�Q����0�|�)ՆV��Y,���I|ַ��3�Cy��#���o��)諿e��m�| �6��{��DpN>��Q.�G�+�>b�B�s��Kr��ɵ�6u�su�-�	߾J<=_Nb�Db��U�9�خ��3���X�<&����>Ի��w10c�HDI�0�L=�-�v<#"���)RkjJx��y����9�����"m$��l���:Iw����5~�����`��\l����!{=�ٟ�8�n\`s�-�Qԍ�E���ބ��@�VB�_�S�Q���8���h�0Q�I���%NXY�U�(y-_�̱�!{���{8��ja٣@ꔌO������X���b�0#0��	b	��n����2Li,�"8�_��e���mn��^<>�ZvY��T�ȅF��3-;�[�^�i>���i�t ��X�7�z-舱a`b��ɖ���#��"g��&��E	�H-���vC�.?@�2�K;ƿ:��]ܻ���[4�+�f�,�e�y��V'���c/ْ�x�U#7�1�/U3��mGG�*��a���1×��˘s��_ppǿ�
��I+��}���`���-�6j(d�c��f��f���v'��ۇ�<2�5|,��y��a�>Ҡ����?(�T�o�3��G�b�y�Z�-}��8F��[�@n@����Q�[I���oE������ť��sww��!�7Q�I?I��=)jʱ���,�Fˍ6STp���ƹr�-��濊�O,@'��Ѷ4�	 ���u>Z�/��L���aknٚ�P���E�����Z<�l]N'q�dYaV>�$�-�e���B��Oό�*3>"Q��C���g~�І�z��K�j?������x#E�O����9xL�c9��ŒC�G����\ə�W�Zyc��w�rB^�tQ �-m�
����fOv��Z�X
�NtG�ªlj�$�Zp����T4�=]4��I��X�9���K�L\�#/e��ӻ��k!=��V�@1�)E�F&�9`��¨�	������]��>e��|�aYy�bKyӓ��n���1A��W�#�Q�w����~J`�+�I��C?Mk;���[�=k��z7
��O��s/g���b���O�ʦ:��Ƹ�$V<![�Pb�F�i����޺f�=s�
���4"�8�~t��-G5d���,���%�[�~��E��ā�i2z����i�h ߲f��wT/�uŪI�o�}���,}�+�_[�*�l�b?Y�~I^!�0�R>��\��2:�gb��-��(�ѕ9j�;ms���&�)_\�}Zr(�����]VM�������y桵�U��h^=�"9Dk�u�d���㩜���eD.9$�b��O9�R� �׭w�-6�DDL|�Dnin͊�Ra��y��-j��n����J�A����9.9�����N�F=S�����ҙ56a��4.v(��K���S���d��˴-�W@����d�5������Q��	q[��2k��]��)*0��W��t`q�7F�c�T�44�u���k.�@|/P� *�T<���g�[w�L7��ztU���^�u��tNSٓWђ��}�td1
=�������7K��Xz�_HpuKx�eB1e�I�ǈmbH�.w��R<#��ya|�� ?��[̰�^�X�
�^�_j�N�����x�N�b�)�T�nlq\L'���_i�F�qh'ZF��Kֶi��k֭�=IFk���*�	���T�?�q��#ѭ��ųuMzh��}U^��w��j?_��|�PG��X0��"�ɲ������*�����]��+N;��#����r��ԙ�D���(Pg��.~D�p�F]»h�q��_��{l���m���8?�aj�r)��"%e9��
���qlO(�֛���+�ء�`2}2���V4��:�́�@�F�i��;�T�>�M$�:S%�)}�J¿��4�y^���va��nN��йF�ψ�4��^q]�4��rP	`�~��5�����+�\�u!��Dz�?�x�	E�N��H>�H�dAO��˯ ng��wpɂ�l�
����wSv����8��Z3AG]���U��>�X�v��2`A=죽^������
�vQh�Y�G)��7E.����P#C����ZI��h��f��2_��T>�r�e�㏺�����W8���H��T|�Z��;������ջ�N#a0��6��I*� 5Ho#qn{Q�,��B�+�>�v��]efY�N5ڤ;���1���. j���$+H�QpF7<�SH�9�D��7�C������ 8��د/����NJ[����~�C���gG&*������G���K� 1ɀ_��m��,ZƝ�b��U�*r�r�PL:<�O�}��Z>�B���>�$X�gT�^�=AR)���~�Z���uF�T���)<�<H$4��#�"�FYZ�c<|xܽ"4h@�~N���E�`�x+g�X�5D[j���]�Of��|�-�M�ʷT���n"�܎>��"Rs���)4�1���Һ훧Y���Z����P���#��2�	��:�Lde5�ϵÄdm���x�S?8?���#�5����3��3��*�ĮdFc'��e��oZf*�.*��Oh�l�C�1i����$P�mpQ���=B�SƯ�k7�ε�]�L|}�˝0k��1��M&lI��du��Pp_5z8@<��o爍E����ʟ�U‘h}掬R�}�UCĩM�z��|�� �3o���3á�v�.H�� _���NUf����B��ʵ�B����%?2F�H���Y\=c&l���X�ٌV�-�Nx����+b,%��9z���1�VO�#��u�������?(��o�/���C�0ckK6�@*��a�rR��'�A���� ��z�+�]u����'���Lu0���B����NmA�����qpÕR�����K���q�[TO�Y�"�S����.t*�t=(T�Z���Y`�~�ِ|R)k��l�*k|���p�RU���)}�2�ը������^ZS'˓��BW��Q��O.a��?��^�Xd��QXk�32lv!���i�ߗ�L��dW$Y�2��#d4)����E�*��ݝ�S>�\��~�	D�5��5��$ � ��h�݆��F)����m
�D��-0�'�T�{�~'���v��(�#��%SэW�:d��'@�x:�n���.p9��7��X]��F�v�򕖝�c�h�=.=�:Su�� >ca�}ѮW� ��*E��y���0Si!#�g`{:��c�]`��mnI�S�l�47�{�4w�� k$?a�4]�����+�c�GKg�wlA���� "�"��SqKz����SY�a�n���j�9�8��ъY� ��_��`5��-.*��`��@y&o�o6�Y١`���6�3�f���bR�����v���{R�k��HZdE�ٰ(ɧ����9�hhY�>�E��8�>wq 󩠧�D��� =�W�l�8� H�9h��6��F!��`V�
p�3J�������+p7�,0�������,W-kZ���e<�r2l�n��gZ!�������c\�;l�Z�`�V��e��v�0�g���!F����d'�N{�?����1L�gC> �I���H`�E�m��C3up,Qչ*^t=v���p�:k�\�*.��{~����[��q���0?��\eN욌���vUq_��Ρ,�8ũܦ��%�j`����ts�|�0�6�K�x=�*H���K���T�X������'+`p������	,dU^ O�j�wv�-x8�e �%c��f�+�����_�:M��t���A*��י��u}"�|a���-|l��Öj�
�����0����B�7RV��^}ӡI�ڨ^A��������]B�`
@�2[H/��l������Y>B_��*j�*�A���{�^;�l�u	7�L<g��,��;���Q?�t*�C��z������[8@u7�]�2�f�n�P��p�x�:W赯�Z3��,,�-���w��.�؟fC�2�?���.u�	�$0�o�/���ǿSo%�	��1��2s���u��}mm��T?d6���aQ;��ؖ�<�c!���Y[4����j�o���mjZ'�A�2^�5�w���n|���|��
:��pul�Z��Q����N�"��Ҟ$=�� G	|��*6�]������-}�=M�PVA��$\����� Y�vۛ�	y
���ě�L��J�k0޵�՟�,�������l�IE���;릹cz\I�<=���sM�}u��Pbx}.�,N���z=*���ƅ M�'�l�'z+*?���Q�;�q�Z��(/����� �} ��A��Ҙ0:Vg
�wf�q�d�*O�0�#�ವ\��X�\u�%.D�fs�լ˥i��?<��]M�V�"�,�Bx�9��	^�{���;�������#WOTy%���X���j�~�y�5�p��/�N�clZ	=�:DKm�8��k�;&5�SN���Þ������}�3�Ӄ!�2��EF�0��#Ë����.��R8.m\�3 t�����~�7�_pD��O��݁@�t-ǚ��:�{�'I'�,E���\^u�q+�F���d�1~d�:�"��]�7�̖5�yY4\�I����鹪�w#A~WE��.fm���)��j}Y]�.	�P����h��T��U<�� �7{h�n�e�$vԶ���h�����ڏV����B�7���h��?��@�;/��x�:�kjw��@K6�u��៌�UNk�l�O��	�q �1�-�Pا���,��8�ר��4
��=�F�b��l����dq���$m���c��.k������H�����q8���bWir��ü-��˘� �z���ZC�"���8U!���o3�kH)��3�j-^\�Kσ��� ����b�0|oO���C�����#��̣��4�;�\3�� �5m��ZT~�?ͩ�]�4�8���Li���B*�0�#���u�e*hǜ�9^Z�ۂ���qAR�'#J�IJ����5�wGj�m ������5d�»�$2 6��w�4�'�� ��t���ō}�T[%p��������4���#N�E*�4
�+%�L����x߳š	��v�XUtA�bi�t����=�xk�G���-H9�j7Е*,�}��=�Ɏ�m#NGl@�ׅ��n�ɲ��zمk��=C���?�ӷOؿF�q+N Y��	yyI�!qA<;�[�|�cu�"I�D��-�p�]ղ$���H��xt�'�j6��Wa^�B]��@����6՞�K�1�J.����LC�dN��ϭ��t�vc�}wC�ФI�l��\���2`u��H�79F�?�l�T�1P��5�f�t#�)�K������H߇MQ��[���<�V�Pv��=�w%�	�6r2
2�[96���ѐ��|��E���O�
C2��G{�-�Z8���5�{'RN�ݱf������jG�a��9���N@�O��c*W�����lY�_�&2+4&�:���U/�\�6��+g�����EM}\a�{An?���w5X�����VҞ����6�*?h�y-H�Hm�CVM��2�+>Tڐ/�,L�M_6uz�GG�.�����^��]�'�ł��l����l�ǻ:~O�k����D<S�� u}p8��2���$҂��tQ�UǠn[|�y	s�A�0�W�D08/�&��ch��YD�H��Wo�F�ћs��ݴmj/����-��O�1����cϠ���l$̅PR��?M�1A��9��� 
9>���e�>��H�Cw��Yw�p`h	�]W��/��4�o��G@)$5\@T$��f����9��)�<G>v�*Z�w�p�2q�N�,ے���7�X*��� $���)���n.d�M�l���8�(��)^S����Iצ�"���M|R39������ԔTΏ���ƅSla]�)�^�>Q�%,�сVXܡ�+`����R=�� � �s�W$��h�[3��ڶ�.���W�ܚ;��Qz ;�Z����.vթ	kq�"�����K��:L�
�%�쀘�v����JP�ӣ�Ή�^��u�X�Y�깩ѹi�.QfK��9�w�*'8Kl�Ю�,P~8��WqY�� a^i=�W�}4WyY?�}б�*MʍGr+]3��O���R����d���\ה^86��괦*���檺Y$:�pF5��Z��V-p;T� ���\���ԙ��"�8HP<�j|���`�"?��e��+�#;�
	�E!߰���If�ccP�1mq�������ʯ5x�*�,�����.��Q]�����R�Q,��W���u��w���zQ�m��l����Ijz��Oy����|B�8)��#� 8����"R� 
���.�"�t�F]0���=�,��TƋ��&�����Bt*����!듃1�Y���<��]MƉ[��q�r��D�cև��t�67U�#�`]uE�>o��#tT�u%{�=�Qh�מ�W��M�J����)TA��خ�s4Ӭ<B�c�v3��ܽJ���1�Y�y'<�uD��B����0
Er��^$�=j�" N������9���d���<�%vJ�}\��U=�9E:���JUĘh�⺎�hd�M ����Jq�3��M�ۜ�'s��z����`�QSU0,!�yo1�T?$Q` ��N����%u�(��b��5/��X	�R
�F�3P�w8�y����]�����L���ަ{��&��(���#�/�)X��R���[�-���s�i<j9�������܍ɪ��Sn�������!J����?)��	�wCˈ������կ���C�6@���@tLK������<�����.���C������E o˹5���3)��x'�8��f`��Mr��\b{(�źe������' �Ia��Ȕ.7��pHr��a�8u�G]�7(�=2;P�ii�]`��9fCy(D�/�����/��~r��B ۀ	y��""�X.���νKIG=J���D��+�w�)�-����y����ǩ#�?��6.���
gp�h��f��CY7�+��">�e����U�G�A�����2��u��7h-����mUexTQ�� �Q���e��9�H��87f��X3ZO}bpw(��g_��;7v繝G��\�R�!��<ӺqÞ u7vo���g�z�6��| ���{:U��	�����j���}��;�=�+{	��WEEf"N�:��\�e��V���.�CKj�A��P[e����1_���W�Nb�zJ��,=uҁ3^c���}��7�3����Ȝޟ�XWC���	�̱���dҟn�7q)�56 :�Һ�>���F���sJ��8��J��j��WnK�b��������$#�V�8H�mbbz��V!4ur=Yj[wRϾ7�z��j����.9�)��.��f�!'g&�������Ii:h���>���
y�(�P��KU9���@�o��9�=�r2���V�P�z쪊�	�!r(
���p���F{x��	���NOH�ϞBflh]\B�a�7��Z8=�>Л~g	�uvm�$ґ�Z�ҪL���7��%��U/E�̲-�^�CUbV���<�9�O��s`фg�Q��˵�{H�[x�glp��R�����i�^p�IUB�(=�<��z���L�) ����7�@ô^al�_�>}%+)�L���(9�Te�Z��e��l�0���x�C+7U��kRp�=�dp*QTF`��50{[��(�dqNͲ��$z*v�G(����ic=�o	���4��81�`1k����V�b$��!N���>���4�q��ZMlFm˙b�N?Pݝ��,Yp��@~j��G�lUť*����A��زδ==F�#��Y9�]�	ݼp)��ep�9�ޏ|6x���(6h�Wiܟ��Й��w.�
���<���� ���Hh��s��*yi���?K�����㋞�ՀR?h�d�y��x0<�!�c�h3�� W������!qS�[�I�����	�O��ӣ���7��\�)��XI�sWȍ�}�S��}��������A��Y�u�`�2����C�lMגy,���1G�9�۾��$�je��40�c�.�گbRN��o;lR[�D����͎�/G���'�� �D���RrL�;�d���[䝪Z��g�<ldL�zG���+?r�6���y�0Ww	!���T�'����Xxg�G�7Y�A��`^I< +R��S}����8�o,`?�]B�F�B�
Հ�UН3b4��&��{lF�l�3ųMؠI�+�g��p���f�XSȰO嘅��§&�-�!�	��sg�k�5+$SH�Cn��W��ֹ�V���f�F!W�y�e�^Kܼ� 8[�J,����ZUr��Z"d
��et���wD/�b� �rw%����]qm{��`���_VЬ�O��ܮ�S��(�_�WuQgy�0bK2e��{��/�@��6�����=��(��3{��q��A\�ZLT�~�E1S-cE�a��YsiO�k�^%���d:��T�%�bu�ʣ �Y�4���@�,_����f�t^�f���A���r/��r��4`�����*3(�dXyĠ��-�O11{�܎�޽������2��g5��h�	�r�-m���j+��v� ��o�A }?�5��Ɉ3{I�7���$PTm����K�e���l(��B@�x>��u�-��8�a\��=OnQξp f=Yt�v��I��EZ2�G�~nm�����sH/���~K#�e��M��&;�Uz]�\�B@IlB����c�}�ȫ4��QԥwpAS�m���w��Ol��P��"c�`��Y��B�Fd�9jp��X~�S���o
bZeX�K���}+��^�RSJ�xU��ߺUx���a�鬅͉N�|~���>��o<�=(���ؘ>��Ih��FYsX%�[�k:⃾�)��Kݒ��+�sTLW����Yp8�&��8Ѹ'e/g�<�~�$��o��{�f�l%�	��5��	�T�:^�F6K����RU-�|��Y&%�П��&���̦'P��� :J��<*��d��#%�y^ڒ����Pm��N�TrA;d�z��'��:�8�OW3�ӕ%�)냬�dX�?����o�\@�r��3WU�C�'>���ܳ��zP����(M ؊T��bJ9]�:4ȏ,	R��(v�l�w�U����[BSP����i�)�&�[��M���V,�ٻpO� ]�d�A�
�>8���s����^�����J��0�:ˬ��JrPYS3�\ug�5^��|v<'���x������m8V�]ie����SĨ�L�%cU���J��c�Y�Nl��f�����I����*�c�p�����}R߸H2
�+�Y��4U�vX�'�Y2��B��[s��6��~���ѭ-g��L�U:�L���]"ׯ3�P�+M�8r���kQ�9LT�X���UU��8[G�^��]>��c�{�7kq?��� R��xbu
�Kjm�bkE�61�7�����e�y�@jl����{�7`�҉��M��]ԡ��P�)Yq�J1{`��z馽r��[���H�@N�ѿz�-~b<�3���ɭ�aG�R~1�	�1��v�Zs�$���=��o-��L�D>\;�=X�J�b�ΰRAdo��*��ƣt��v�4J�>Q4߿d�sx�Ozr�z_�noCs�R��,*��K�">/NE(і�9������DI�"��]Ʀ� ��f�EwEd �UO��Uk����&[>�ݧv��PJJ��P��j;�}-Gs+�ʳ���3�)����`��^�z��]�Y�W������&�q���3yV��vSQ���ڟ_ξ�#ZS��+�H�P�̲H��]wȹՆ9�ÙWv�C	TV����_�rٮ�)���[`NNίe����5��5�t��f쎤�W�4e�����w�,q�W�'�� ��Ӗ�C�_8���r�滮?w��g�-��s��[y��{���Ǝ5��<i�+%����0@{�j@�1� ̇�U?�q϶�G;:��jS�����D�~9o�`T�D�������$���~	ٷ������/�Պߖ�%h����ׂ���͆�xkC��2%i��b�i����GO��\�`wC �J�"�9#�渥o�T|ǵ.�pp喀֙�j{ѐR�NT��P����t]%d�vĕy(��h�>��O8!���(��z����~�K����=�ĸ����U�2;r�X~�0Sj���z%���P��wjW��͖�2�b֚�8�-̞Z̩�)��$g�wEv0|��)Ox�����c~"8=�؄�=3-�П�!�i���?���$y$N��Ua�)[�� '��Ϛo9B�����@��j��'�e�٫9�Ў�C
+��o��!���L�G��{`�:|M"〉�sO���3��G�rI₝�(��m�P��|��0�a����;m��`�{�!_�[�/j���uM�@���7<:��~��̀NN�OѨw���egG�+W,�{OLA{�Y�F&VDHG�cH棒�+E���������_hI��#Ԁ���S�����3��+|�l'y���p��T�]P�!RE�t�����QUi��B{�!u�3�[��<����7z��c&��w��mԳ��N��);־Q��D��Ao�B�C=�7`DE�}�e"��r!.�s�A�,�"�"ۑ�!VU"�;pJ+x/�KR�|�;f���L���j��޺b9��g&��W�����E��C�g$ب@սݽ	G���m,�r0E�*Xyq���v�7o2�H����A�Zf�M����<6�  ��3�ωvz�W]@���.Ĩ<�U{ʿ����I^��W�K���Dy���M� �~+�M�W�1�qi�o?��[�m�U7�5�=��
H��t*y�m- ��ջ�B"V�k��ȉ�Q�N�2B�3"f���?fx��Ԅ���hۦݺ�`�Ro�Ϫ����dە���d���_�M'�(��S���r����02��+gvx�gʆ����d��I7�P��U�/,s�oS�
h�*�4�6K�*��Kz`��@���e��;-w���ۦ�#	t��mi��)���t)T�i�T�G3��*aA_���n�uoF�%���=4@n�����9��6���� T]��)��"�rܿҞ��ݫ�5������MF" #x���ݗ\܄�Yϫyb��yC��߉sO�[�6�8��TO��t)��&�R�T�'�_C���|^K*{k+���e��������
B�q2";U�q���Z�Se�z��Ϛ��:����|~���3bg�<2��(	J������=]�iĊQ~���E�hN!�h�k����^�_��>�"|N~���R�|W2�ʟ�X��xvC��?�^TC��Q�\�6#�Պ�g<��#s%�N��.�>�MnAĎYf6���h�(���:8ξ[@p$�.� ����#�'#�+�X`,^:{�`�d��y�E���N��[��5"9�P�G�٨�9\���%3�;��	\m�]p"A+����_h�CI;��?��5׻I}���IJM8�K��?Vcᤆx𚱓l�k�_�Y�����b�0F-�Q�kvQ\B�G�n?�0%�K3��Ѫ�h����m��8'�wM��^ע����XC�c���3�j�͓""��(�3$WE�>UƜvf�s[ֹ��Y���)�/�_�RR۷�^�0֡՟�O�����!���~ K�-�(�� U�28�^�PZ������Z�
4�X��9w��h,��<�@|tI7:�Q\���A�v����D��y�������JJ�*���*��d6]���� >�٢�?5`�İHXB�K��#ue�ynӄ�{@��i����,�\��ڛ��F��4[х7^}x�Y�O~[/m�m.�/����&=0N���huG���.��U��Ώb��'�K���l�%�Fޑ;������[�&N�j��@��/���ga��R��ɾ&tF>Z��E3���$�:>:�
�to�3W���B��,���1(7��"��s��[M舝��hv�[�p6�j%pX��W! Y��ht�2õ�埰���������K΄���$ˏ����B#����Bk�6O]-ƙ􉲞�r&g�s�3�
{�H��L����s6�nE���Y�̂�azF �EgX�3���B���K�L���wG��1TԳ�x<�>�w܃������f�b���9'a�+��y�ׂ":�UԫJռ��,��zmP��t-<����ׯ�au��Q���+�}˶؉����*\�g5�����|{j�Jk��]�'EzU��^櫹��g�����pm�P���}W��@�=,���B��	Da%����?�٬��;�8�A֭B�0�.-RT�V���Q�&)\4ؙ��WO{��G�u��%�)+l���а�Dy÷W�����ښBK�Y�l��N� � �+����'el#�g���^>I�ZH
�b��*hk��C#�u�k#S�V>����bo6Fݬz�ѭ��������%JH�6�ڣ!�@x��z4|�v�葍��:&���GC�+�6@.*���;ժ���_f��e)�k�M�8��P�BǨO]�B��,J ��01�:e$�Ʀ�t����W9��a~#�f�vB�//?��S"��5F��]��w|˞�k)C�f�#0ް)��tG<8}Z"���%�٤I��G�^X�������܀T���}���
��j�$F�8]{����l%W�(L_Oi�YYנ6�;_�0jǹ7j���U�{����u�8C��nK�kt�'1
1N��.�B�da���޻�����¥ګr�;�r����♰R�7�Rā���U�Q4��W�Ė�ud6z��Ē��	�k��%�=Qu>���
5�4�=3���c�ѥ+�ſ�`�������:�ԑs�
�I�ݢa�eP[���S�Ic,_6%��Qu���e��i<�F��j�|���+�Oe��LT��.��`!��Y eَ��6�SG�U�Y>����ҜUbx	����*�
B1s��n��薭���eR��E\��bz��U(�ǻ8�����gE茺��8��'���\D�K���d�#r�H�v<� 	\[=��C �I�J=׳����]lvv>��dN�s���Ƈ,d�xr����n��	4�������fqG��#�-j{�V�h�;K�t�+	`0�ލnx�&��������
�ki��r%T���e�	�ٝ����L�q���kb�-�D��{�a�Ŗ]�Q�lŪ���aLKh�U�3��/�y��VS����y��M*���?����]�����SLJ�b�2j���[��T��L�:8L]r�g������Td0�����UwB�q��MGJH2i
�� ch��%}d�a���"�@!^�A�P���Vk�'!{o��y]���	e��}{�|���H�R.=
ٶ�x`Ú��hk�Ru�-=���,x'\�`���t���wE� 1W'����<&�:,������uj���:�H��8�?�<�X��m$���@��5 @a@-[X-o�V�Waf�S�e9�]�+�|8�N��e�%���Gn�쳳9���}@�RmknȢ�e]H����6X�ͪv����n�c6
�ʠTM���b0q{a��{/�&�5v1� ���l9f�a����=c�R�N����A:|��ʗ��L�\�o��g��U�Eۣ-���2���s�U�3="33��v����=���~_;O@ƈU��y���$�	�I�t��ZхJl��J�#��F|�+��bI�i�}r�4�B],��4����-�j!��>�~�La�k�o��g��W/�#"%�U�k�Bʰ�����o��F�O��L<�}
A������d�(�X�=P�I1�v��W��Nd?!�,�:�U6�X�	̸�I��+��wM�=Q�ݥٛ����sg���E�=)���Q���2vΥn�cTN^�6o�����4����jC�"�ޤȫ(�b���Ȥo5��W�$��������mS�I� � NU�2�ݹ��˦}���GwE�|�P�ab�C����CD�M?�N#0������oZ��:n�&7�y��!ڢA����/ d�b��Ю�R��ѝ�Y/�ݩ��Kȅ�c7�Вޤ���	b�XE�t4��W.��჋VCC����Z73��t�R�j�"�MP�Z�q���v�=�$#�"��b�)c���>�����Zm�n����q�����|𵆑@��nr:[��f��%������N�Y8���@���"�ϻ�E?D�cC���o���
�SɭdrI�^�,��$�ש�ʺ�8�;	)�kܥw�-WkQΰ|h�E5��Ps�O��Қ�s�$�o��TOSE��ia2���N8��=w�6�(i(�H4�E��	���HG�#�{�1�}J��=v�I�fs�vH�u9�G���ȏ�I��b��g�+<�q��&�8��MأV7~'k}b��!y��4W����(<x��K��-l�H\���u��9]@�hT���{�������ed�1�YZ0���l���)�!�Ƿ�t�~��jo8`'j9�#"S��}�e���0a��H 7����u�+�D��[˶ �컡�sA1f˩(:G�#}s<�A2�U���}�_"�V�$`��hN�?��d@� X��dT��B
�נ����Q]�:�V5�~TQ	1Z���ohc������I@�|�`Ӕ��N�����^�-���2�?>�(�HR��0��l��A���Nx�T��J�;��`��oߋ�5(�jTG��j&�S���4)>����7�����z�-cȭ��;v#����R��2��)� L1�%>U��l]lgq�a��c*����r� �Ls����k��z^mAG��r8ƭj�0�H��E���	��7��+�c�	��}�j�.;9K�F9�qp�2�Nf���Tg��|&'7uA�ᩒp����`�$�"��U��i���5<w"͍�%9�}Ǩdd;"&��ǧ�ꏆڣ�c���þ��&����s�߂���]�3|/�dHmhzod���}sg�_#��.��!o}�!�>����^,\9��2u�,o�ѕ�U�� )��o���L��p,լcWD���ξd�y��B�.{~�r�)��fAKt���� �^��Y��Q�h�+�|�א�Ù��+6�]�f"0�$"!�KnC>$_A���}��-a����ų[�^�m3D��Йk�`�'y��H^��^�x��v|%e2��iSI���0����A�!�J�M;ʤj&�Fg��u'��
m�+�����-�lF�$P��C;ӝ��%�h��T�$��mV9M9�=����h�m�4@���e& ��YT����c�Jy����x���_��~��_��̉�&���Yy<�H����/��9`�W0���5�	c��iB�ə�A���k�(Ȅj�i����T�� ���p�{��@��M7̐�K=mo�f0�0��)�~�anrGy���6�~�R�D��b��,��{s����0��.�p�� ����u�����"�{�e��.t��gI�z����ŋ��(���Q�N-���)jS�a��uw�T�&�8r�9�ͪb<�Ez�e�`1Bǥ�;�u�q [��Ld����0>��+��&%���I�d;���nb��RM%�[��p���of-��v��h0I�bl�t�����թI����}��D��Ġ�y�A��B�W���Y�ogo2�^� ��V��xP&km��X����E��a6�1�|�o�M��A���ϒ�����x����vVc�V��T���o�v���H+������3#�9��}��{��k!�F���ȡ(�u��1n��C7�|����GA9!�aa���}�H�顯�h2�@���av�v,7�r�o&��Jo] v�CZ�P�\=�qȹ�'�V���YQ#�(@\J$�>s�.�[l�{l2���Ӱ9T:"�x�EbS�bgؚ's_?�B�*m2�IS�p��'�@��x>{!�F�rk���=��İ�淲�.�i;�%
�n��X���}>�=0���#���5"��F�ǹ�L�K�D+�
���4Z�,��C�Y�T��vG����Q��2��,�Dm!Dz���Y��q`� �^����r��<&V�?��	�� �+;�!�3@�4���ǚ�m�v@7��ݪ?���"�z� �1"!8�Dѷ��t����ģ��U�� �v[X����m�?�_�gan�t�G�<��6��a��_�o9\T�洺��:U����f��1�ܠ�
q^���u��3\xʤ�=���IĔ���b=�w#硠>��Vi�p�l
N+[����
��$��0Fٴ��$��.�C�$�$�����h�fN����\!䥰��Aȃ�9�5�B���A��x��.d �	���?B��UCK�l�߫E7I��|KK��D�q_���Y-%���ec��[��;p�#M�h����T�=�^�9Ճ�{�Wb���bI�d�}��m�8��Ea�)J!!찮R�`N�_9�Ƕ	�o+Z)�D��~M?&5*�
���%�>.��w��˻�ݳ:��l��:�ɜ!�����#�B$�����P2�
4]��~X�%{��j��J�<ȭPC{<l������
(����m���ݿGE {����l��`���zҔ���6�|�f�s�B3���(y'���bG��ڨ:������=�7hDm�沙�Kxz������$ J�{�®�[<�PLe�����#�.[��ݓIJ��S�`R���2i��ch���;@~w�VP��jD��{M��e�Ԫ\���_����Ʒ��i0H�a__�nUL��6�n
�L�p���=&��wRz� R�t�A#d7D��z�Q��RGP�$vs��6��g=O\�i!���D�{���H�g�Y����X�>ˮ��[`j�н9@E=�쭲Ƚ��,��ޣ���E% �jw����R��(��QpM��=A|�\�g`��9c�cß�X����
lcG�<`!��j	;&}v��,L���l��3Z�}��hS�C�7���HZ��V�v��a�������nj�*��=�-F���Ac;�n�\F�׬�K�'*��Y����#TH�yCǮ�[@gPrOd)������G��A4ݾ�M���y��(�H��v�������m6�_4��v'�o���.�8��OO��,+g��2����s���M0��v�" {!��I?��3�y�Bk�YΓ�nt7�%��V�	ť"CVH<hh�L~���Z���\��'@���2��`��fW�C�&E�.�DV�>���A�0��Âdy�08��xZ����k�Y��|����+6	��H�?Ŏ��u��L�J��qc�Uq�P#��&���&t��-v×�����5�B�t����J���w]���G���R(�;��gǰ3��=P�K�f�@���>�y�8d�����g�n�Χ���'������VW���~�	�Mr�L Z�)F;{|��^ћ����,��fc��'��yV��U�-�r��/a�N����|��f�|3�V��Hђ�2�B�N[����2.3l�-h�kY�^ ]���-[�U'w#$�TE?ldgTH�K��� �1^Rp�X�/�]*w5Gl="���Lj�0}5ns�Z�K������]d�e>!	�A'p=���9��+��1�$"Me2�>�&<L 5�'4�BɄ����ZW�}�Sk��`>��RH�6����l�HoL�l�(H��[��
���W��3�w\d4��#3�4U��ƀbsi��\]�ZI.=�u�a�L�W�������	�4ֺB�q6�OU�
��tL���3��w^?O2\��0�,r������S*�`��?(�<�T�mC�p�@0��eb�_�B��3+6 ��eZ=���Tlx^��D��v�4z�6,Dފ��QH0�ʌ��l������0�-�KfiF�b��w���>��]�I�B����rķwK;�����m�i�KD�I�o@������z���J���@R�q�23��)� c{f {�Il����
�����������+�戩�����WK}U��p��π�BV�f��$��o��Ci��cl��(��! ���oիks��EAw(h�SyJ�G�X��������D%�����ܓ�����NX|�w	����ś@�cl<�KH	ż�nu^����<�x��Wk�LBt�����|"a�]���t���W�����+�^�JU�\����'/��Y��@�
�M�S��8f�����00<��FުEǿU��h[���V�q ��%Fm|�j���==ٺ������il��a�M5�2�uHs�b,{>�+�Jᤷ�j�z%0���tS�OXQ3[������J߅�諝dlpE�d�]r�郖�����	_�6����mcf[Wc��UM�)L��q,Ȅ��>��t�j����/e^��E��2�)������w��ޟ�J�=���a~�������z�Uֺ��I�U��s�k�[��igj�r�(��'��5%�4#�^QJ�]��?cB�Ki�B?��@���GǦƦB��l��)L���H{��e����c����;,g 2(X��B��ǡs�9�ޢv���}8R)m>C�����A���.0����E�Keǿ*<��s�#����t�p��t��{�h������� �У]��-��jp|�Y��Ei\���Q���a����at��Z���>�6R���6d.�L��]Ĥ��PqG�%����u#�=g*><
SA��s��=LH� �ퟝ[[o<�eA:6�ٵ=���Ӂ~V�D�Q��o �$���)!.P��K�s�����ǎ �e�Cog�r�,�䴨�~�1�',�Ȃ�����?%���4Q�{]�a��k]�y�����N8�������*�V��u��p�%��6�Y��g�Wpħ����eU�5~ݻi=?�[0��+k��n�12rՑ�"���4!Z�OL�����tf��U���J@������� C/�& OXl����G���C���r���"��l;����O���J�׽㲴{�F��t��o���C�r��U��U:�ȸN��e�4h�q��O/����G2�i>���	?���#s��IW�OH�n����Jf	O7�o��!c`�D$��~eU0�r"�H��g���P!��_�w��-�	c���0���͋Z'��#b�W�"Nx�`��ot���2B�8�ͨZ��>�yBO%���v�9���I�; 3��V��p�6��{G�r�1@��s@O9)G%�'$w�B&�n[)�'�m�a#yM���G���Y;��z���(l�y�UH�n���� ?r�YCN���x<��&�Ux���Wt[,�h����g���)<Y{a��Pj�W�Ƨ���U�qUʀ�7�>��7�Θ&�UOs~�̍�_��������{X���g�_�A�e�M�h9��.������IĲ�uٜ���wyzJ�zN�nj�2�o�6xj��1z6wђ��Z�t�&NǊ ��z1��Q��B�j`ԣN.W�TӍ^�.�9� ����ދ�o���"w�I���^�L��I@�P����":����=���K���ƚ=]�X|-I���Kr�b�v�~<� 6�Cp�.��Z.;aT/�_ B��}a�E=���0��	ׯ�o�T's�q��O�������0�@���\QgP�}�l�X�q:	�`ӵ���(��`E��X�;[��<�����{��{Tûd�Wf]ڹ��;�!�o/<3���>=A������3�|Cc�g�,0
�ǳ���Z;G����o%�N�]��u�����Hg��I� :�nf�SH�g�#����_��rG��!~�~��� �O��nFKX��/��i��8=��n���!�X��B���X��x�4)2����#
�&��z&�|<+��#�N�2fҷL�.��oE�b���$��4s�AH�u�Vj���4Qj=k���Y?���k%�gE+�����
=�e���6e+((���x>���"L<c�-����vn�|�UQMA��J��L��AH�},WJ�2�D��ԣ	{Z�TZ^\�Gn��v.��v3$��m����5��o�,�H�߻zXUc�;bt���u�i�E��G|�U���0��sa��o�Y[n\����(�*Ey��)�<�u��7_�~����R� � ʱxR� � ��k��B���R{Β�9�=�ȿ�\2ڒxwzǔ�Ãv��2C���}��\��_��5�ol�n6��FtP�9)h�#�i�W�c�Ì�4P�lr~��ӼJ���12}�������2����6���bH��O'=EJ��v�T��鱗�>!�~<Ya��Y�hA>�w��:�(�X���	8B'�7#�4��P�t~�<�=��!<����wS�����DR��ܐ	���|��|�����]ʒ���*5�_~��W��aU`�`�8Ч�h��5D�������ǈq���r���l�m����Ǔb��u�xb
��Ѹ�98��C���6��^�ٲ���ecUlU�����^����pD�0�wz�9�(ӿ�8��RK�w�{��z�*t�lhZz���}E�+��>����<�"���3���~�F�,	@����W��ΪsA�ե$\�"H��X�h�wѕx@����� ��SF�ZLq<ਨ�!���0SM� �����H�����Zj
⅘i$H�H~�m�7[�kY�}Q8X&����6�ѳ����֝���.	��9���}�x�2@^ل��.��A�c�:�b"@�Y�V���?��<��Z^v�#p{[5����E�CQ|��/X��vl?�Q��v:GFm�_�=��}+Oy�ы���ѬO�хw�����[�I���%�e�$Q �2O�g*^��r��;�0�6P�Buo���j�v� �e���П�;��Rqc�%������ܛ�4#���wh�"��K�9+�a��c�!�p���*���gQ�3�A��y��o���+�,�E��	�l�*�]9Q�����$�"�����̭p�ԭ.�8����}L|*�H(.���a�Z>���E6�H�Ϭ�w�jM��.�jQ�Ah��9� ���Z��:�ꭖ˺�O�v��+Ew
&u5@�Qܫ��UrsWD��w����UM �
�t�O�;cDB�t�����Fm���^����f�@���E�}�{���`���Dc�w6k��C��h\9���{��䧉���#O�>���hd
��竏t��|z�0`yoϣ�A�rX�PIFX�B�����4E�(��,[Ι�x�`���
���l1B�O��'�!�M^^"�v[����Ok��cncْd�J���tlwU��<����ǋ-��h��'���.�`j��k�6��~�N��8�?G���q�� �!F3)Z�1�����,�9���4�O���Ӫ��Q�E֙��[k��6������|����w����/z�b�H-͊M�z(�S��3_�q�M��$���s���m7�eb%���aN��Yi
"���u�К���x&�5�#W���^��tZ�?F��:Y�A(����s�']*Z����������b�H'mq��4 S"��^��xܠZ~8D��0Y�D�_1&��]yN�}��t�#XU�,s�AWϊ�}%�|��(
6tg�{�|=�=�(����6Ջũ�7>O���	���cg�}OHWF���}�6\.�͹��,4�m��S� ���œ��ۣ�xC�H�z+l��\$Փb��Nx�2��'��n˷����.�u��{Fr��,�'�`�ǆzw�_���$�j^���^�tY��uSfs�%#AN��ܢ��������kZ�]V�[��q�i@�RV��K��Q+���w����,�'0Y+�p�YC���P�!֓JI�X~$��Mm�m�����Ho�Z���O��O��JI�̵WZ/-����$\9 ���f[�(-ԇ!ɂ�2%�˱Z�QO�lO�)���lۜ�IB�*�sߦ��@��kq��p'4��Gc�c�q[����k����J`�9��qf�h�Xfߙ�ʯkt/(�HV�J_7H��(��P�?��e�c��έ7��_/w#ִ����H�������7��)���c^~��h��\���~�
L?;�";�"�ƨ�&\_h������,�[�G�GZ(�?)�Q�;6k��j(_�/T)�5�PKA��⽨���`Ʉ}Ȑ�I�������?�h��5� H����D���Ǔ�B5x,���~�Pj�r��-�a���V؄���X]k��%��]�i��=V#�6V�\�h��Oo3�����D˾n�^�o%1t`E՝�ߞ���ҭm���|Ծ�@�$��
�*c,,4u�lsx�
��}�Qg� Ij��X�Xbȑ��~� ��WT�"Q���a�a�d�`�H����(�@�ȔU�0�NE���B�:��m��?"�Nُ��ه~G@��[IY�L�a;�+:i�8_)}_M�{�I^q�����#����;�f���� y���_�A01MO������xu��;�g� �h>�!%|���)�Z�~�
��� �~V�)GM#�F����CB��WN�V�[hU]���|��ФB W`�a��O�96��j�βҝw��.&,w�}��I�k&��@t���5,��.�Ǣ��$�`h�S��xe�u�L�NΓ��
�����`�������ڮ�0j����g�Z��-y��bP��|���a�9����U8���-��LsX��S�����.'��e�F�$V��7�׾�aw�w�}(��O�,����Jf���'�06s�YE8[I|A/�}}J�N�#ٕƹ�i�kDq&�@8�;�#��О�Y[�����ճ�/Y8��\��u�H����b�:/��l��7J���� u��3��i����V�"���j��"����&V�6��p��1�X6������3�} ���F�,��d5O�CA^a;�_i�R��b X�A ?T���
��a'���[^-�FըQ��,ox**�k�yeI�|�.]�w��j�ÚG�,�7E�-^����#�d��A�\�2�;l�if4����|���li��7m��1M�E�w����c����`-����4�����f݌���P����HBqWu>h�lx�&.3w`�Dܚ�7�E��9�����`�����u���פ�e��jC2�Vm����
���,�֟;Y�������.���d��(�!s)��×!_R���X�$R�{���!�����ܥ={i�fÉ)�R?u"8�U���K��d:c��>�����YG*� P�Q��U�����(q�:��]��"�
� �{"��iE/ށF��m��z�l$���ciUј��c�2e�}*c���
���c��_�smnU�r��}i�i�)�ܩ��\���F�i>WU��،~�|��ͅK/��5"�6��v�Ʋ��R�i�k���jfD���=�y�ǟM�>"�Uz4._~��*z��܀l�Zd�4hmz�Zq�Ų�F;��Dɢ,yjo�9�o�W�Ig�iQ۪�6W'�̲�
f��(�G���������2UmH�*������
���2
ڬ\�j�ՠ7���uI�[�����zE��f�+��:���q�A:�iD5"�+�#]u-N��W�G\�6�Sv���S�O"t����[�l�����Nr��XȌb��� �w�ӏ����j��(�"�S_�W�ƛ����9�q���%��t�	�����#�A%DejaȅY)c�h���"���n���Z�W" �Bٿ?�=�D̫��q�����{���V������@�8��$��s�}�ߋ�%e���X�Ҟ�	7�
!�k�����4����O��8F�rOܾ�9�T��*[k �mZ��OT��k��_ɩA�=Ir��zq�2$�@�d"3oS�ڟW���Di�w�6�z��[f���q����
z���BV׿�<lu{��Ű�r�pVǍ�l�󛏹G�B菇B�w�����/��:פ������	�vUժ�6���KT�A�<L��]TcQ b-�4�*�Ej�1j�gb@Bї�^�";9�4MNUHD�#�����C��F�j��	EnF`�����FYR��a̴t�KӠҜ�z�zA����O�����"{���	�����p��-�s��=\�E&��P��O#),,�'�#���A�r�4�8#u��z,D�',KB����~?�4��{��Zs���;��0���3۹^�9��5#�[!����nFbZjf�9t�N4#_�F�TI�Q�9�C5}�ǰ ����:YB�J���^���oE��Hc�h÷+���´�/�ü��IGշ��U�0���4TqE�#"���D=[�����L��oT()�(��{��i�����"��&s�r��c]"�}�US1���`ݧn�ݗ��!���>�.�v�|z��c��OrA�D�E����}�%C�)OE����a0-0����i�q]:#�I�G�q �kk��`��7w��@aT��>�w�7�N���D� B1�T1^�u3�II��x�	������� �r�%����R��W�mf��]���v.#��DC�F�('R�z��Y�.ć��C�Q���:}<�rC)�w����@�9�!��a�c���8��=�L�@Q L��bTk��3���YK���F��y�u�l-R�(J�������sx�!9d�2�dp�K�@n4{�����G���?�2`}t(�F�����x/HYv�*�-��r�;FS.HUR,hr���([]?�����Gn�~���ވI�y���x��P���E�]��<��O'��r��P��7"�3lzϭ:�*>S�*�%�p���{Z���/`lut��<��M5?^��{}ڪ����sUL\���EET�oK�Z��p1���W�1bcW��Ǭ�i^Re	b���?��1�ʺ�L��h��4s$�jCQ�J���|v��t#��^]}��?�����%�R��3w��{=�L4Z|F���I�w>�h\�)C�F��j�f }����I�>�o5$��ߊn�hH=/hC�K
��O!���T텉\�O�&qa;^	d��3M$$S��Yj'���s�-��������R���»Kf�����Q_~@�'I��-�O�i#�*7[^�v�#�kL��Ikԕ�uƎWg�+�����ڋ�q�H�xy����g�YӯG�؄#�/�b�bsd>��<Z�^�I:��-O`�9�yb�䧋�7,�V"�i�G��`-sFY�3:H����mV[}l�9�Jz��Jg���F���/]Mhf�2��
��]w��|3e��K:h G�o�@���GO&��N����2x�֑@���9ҫx�5�P���5�!���5$<!k�͇c(��z-��.�5@���i��Cd�唤��r��q�N�%&�ʦXR��[, �<K���U��Z�Zm>��1F���c;r0�:B}�ʠ[E�^ۨ�Ik΋��^k|��6�o�Lm��0T	Uqp5i���a��������g��s#����]�_�����	)0k���r2���Whn��4?�e��T	&O��$�.�p��s9��l�� ��Q5Es��+Tc��Ik�-�kb��I���J�^n�w���)�zˈ�]��`�?�Q��Q&Pb�Y���s��R߱Xn��ޗR�a�w�2�$�ƞ�^r�H�|S���8�	�%�T��s{�*(�2vu��T)�#����m��+������'y�x%��[30���G��d��"��J�é���)���B->'�sw�OǬ��6��g�WR�@�>���[v��T���`c�z�������+M�����q7�@�#�Q��yV��z��>�+<H�.��>]^��~HR��aɒ>l�qN�Yd�!��ga�G;�32���x{����)��[�̨,p��dR�W�b.����>���$�����Q�	��b�T$Z���}�8����H�X�7�f ����[5y3$���Q���q!�4#��z�����VƂ��=�)�wc[�a���b�O7�h#8��������c�v~-D3\#�3���(�*��Ώ�QAD�Β7tZ��w�rC?�F�\���2��w0�<�%���(@VIF�m3��c���
�B���,���'ヶ׹Fo_��ǌ~�<HBk�M
�l1�1������
�+J�Ke'����J������=W0��l�R�O�(C�{��[=�=݃;LP��v�.,����a63�Ŕ?�y	t�� /�B	�Iyw��.���݃�-�� �b�Cd�L+�	��=r`�WUO���6�0_`����fآ.�y��� �募�wbO�*C  F9�8��;��+�k�;��)z'.���a�}ͮN7{��#!�N���T'��V�Ƀ J���Z�L���
[�2�-�ҷ�_����YJ�< �c� �n1p�1�AK;8?7�h��[��x�&��&�C�%����\���h�z�v�x��#�M+a�,�c𖩊Ts��[Y����r菍Z��7��@���,�YD!��k�����.`�`M<�J5���$3��v0>N.-t2VJ��n�=�l���bA�&/��d��!��@'���/U1TIަ�(��Y�{Ow�f��"]_dw`����f|�Y[���z� ���Y�u(4�죯��O	X�{�ۻԚ�Ω"��F?� ?��w��}�.U�<�7��V	�0�dD�JP?o�*�����AoeW�D��?T T�~s�i!Hf��֎ %x�ߒ�F�=�N�j�=�QT'LE�]�B�[�*֚�������]��0jb�ep��Fb�p�]�
��;����b��`��:'�_�6��ņ	E��x���I/<EÈy�Q�K��E� ڭ�V*�����O9b�`m����"@ӿQ�<����^��u�c ��5�˻,
SJ�3��V0 �S�D�CRS��b���%�|�9O�]�f�N�u���V�����m�q�?!,��T�|�bT^�\����~ �/�y�H��b���a��0D�Ҍ	�-�	C�*����q�H=M!�.ƍ�F��N��k�#/��<
CĨ�d��A�ɷ�`�����y~W+	���%N�\�C��a:�S�!� �1=���ꖊ�'T��rj�����8�ϛ�3B�߱Bݯ� <�3;YQ'��c�N$���� ���Η]Qr
\���cC�=8�[$)�>��]G�M����pr@�M��s�.�,�T�ā �>>�6/WWXE�q呠"��� ��~cd��(j��fr&��Fޫ��a����375�7U��vW�)��E�h�����I��E)�������ˀu��MC=4�O�ĩ�iiF�oKJ��9Z嫅���d���e��:�Z���\���%R�o$ FcPch6B�\���u��XV��膦CE���  �'�X,������2�ܤ�z0)}��(��䬼n����U+������r��=�����p^s̨p��Q�V<(X�"�;mw2���9�s��JEF�Ϊi�6���Oq\M���<ˋQ\�t>�Q��Aw�~��B�'�÷��O�����U*��S��q�#�1����a���묅�t�8S�-�p�ZHbq��GWs�� ��QEr���Ȗ�?�,�-������)x$f� �$ q�Z�;ٺ��kV����������ma0����i`����0�\d��_�h�¼o�:)e;�'����Q��lzNx*N��"�!���J�{�t
���>b� cC�K���I+��хA���h^�siW�_vHrX��i[Mǯ8d�gڊ-���D{Fx�c4�ޛ�Mo�žB<:�:��XK�ֵ��П���ݡ���DfSuU�8t���N�ĚCҾ���\+<�� U�0īǔ XzQ>5�s�%]�K2��cV��LL�� �^�Mo�II���$Hm�:�3͍�h�"�p�'����"�S%x���?I������f�Rq��Ω#��`���o�VP��M�0VY�!��@U�s�X�����Zk�W�~�H�~q�c�#���ª>�Bd��_��nڴ�st�^G'��3Qݸ93S!BD@J�j�.	dͶ��O��1��U��S��IR��'�z�Ǚ9LLi)NN�A��e�-�6iV��C.�	�?�17�F	��+e��9�%#A�R�Z�w��uI��Bp�I��9P%�$J��0ed2[�ت��3~Z�-2me趛��P�&.��F��n$>��~R�ɕ�\����1�-ʒ�4$y!MƤ@T��+��y��.��Hx/��VзI�'�'��7Vrpӏ�+b�~<��-lE��t +��`��v5�{1�c��.1W/G��r(��*�#�đ����L���ON���p��?A�h�jϑ8<�k�S�C�8m�t:����L��(<]W��%�c~��R�O�,���O����Qԕ�jH���ċ�r�<RQV(u6���WQ���ɷ��/}�e���Џ�����
��0���ꪕ8X�'/����'e)�a%��X�s��]�Ow��< U�����qX�h�d�t�ڵ�F�0��rb�y�&��Б�{/�(O�Xm�iX�fY�9,�J�=D�=H 
&o��{�v�n���L�Gs��r�p�H4��S��}{�o]�]�W�S�'é�Փ���ח�v�G�vk#��]邐� �V�">/��vI���,��F��QzhH1���/��(-���ղ!�����(�����!�HR�������5�u5U�m�p�B6�{:�"�O!�/3J��X�R�ZF%K�Nn5����	|H�X���&���&��2���ܔ&���JM�^�@�j�M�p{��/UB���3\��X9GS���ʚb ����V��d��答g����sxn��Z�SS7�һQ(�ꩧ�9�2�W�M�b������&W�k{�����)�L��c�:��qdy��/��Q٩�)7�EBxWy[K�l�4�H-庚�LM!LI��9G�
��78��+��^�Ƿ����r.�z�y�Ǖ#�^k��*cϹ졏 b��:��ꝳ�[�O@�����D�%�1�߸E�i������1F���)�:�+@:���A��13���b:��U0|�BR�����x���Aڹs]�3��c�y q)��hr����q����!�hu6��{�����*;ԩ�f���	"�o�����X����/�0����A�`BP$�e��Eرn}�k�^l�T1�Щ�@�n�:�i�3���JȢ�K��~C�������׳�����T����
��seyb�"�M����M�K���$S��I�)���J�?\��(6����w�wx�V¯=	�����2c�뉷�/V� 7;�@X"�(d݃�&���[�4����it�H�c����b��-O�LJ��� gN��M�*��o�A��Lv��lap�܄t}	�>�
�t�(���x��.I-"��_/*I��"�)�ς�-{�ױeC5uG�*.�����r+�၅),HG����qГdQ�H^��Y ��o���
��)3гy�&�g�X�q�
h���Ș8���6Ƥ+XD�KM�%%L������Gƪ��n�i
�ʿ��i�%�9^����d�f�E�!u���}�y��1��z]n�~�;2��W@�U7���.�+0.�r�N�CQ�|h�c��W��vu��1ݤ��R���s���g�sw4Z����p^\�Y�d#��{q�c-��1,���rmŲ,�p>�6I�>�N������iD�� ��.jҹ!�Z�(��&�e�ҳR�>�g���e�Ƹ�7�bn���\I~r�Q��Du��qǥ���]u(_d$;�E(�����,���{:_�<W�/7�/zeJ�v��u�G4:#Q��� �K�mVh���o��>�����ʦ6��X��ø!������@��%(�y���L�>��tf�yǰ��[��k���0�T�ml|�/��9^�o<�r,����е�K���Bɿu���Y��a�O0����On�.p���]�Y��E0ە�I�>�D��|���߈�.S������\ʶn��vC:LcS��芷҉^9+/�Lo�;�f2̀�2W�R�_y^�����̐к\Жm{�/K���/zNdTL�|��p�ex�2Q7|�d�tH�vokh�}HK���>V7�}���'��ԗ<+/z�=��ם��Z���Y�>Ւ��syTz]���.J6J�ҘAZ���@ u��^�'"�49�����%��m�1�57V�8x)����Rg�k� es*.�j~e��u�ⶓ���/ ���ZDIpe��>�fv|�Cf�׹#��hwF��}OZ�ݐzІ)�k�}�d����Ĺ >2x
?E�T�;!^,�v辩�H�st�2� ;F���`�8n�ϯ�l��U�^ds��UY�?�;t�{9��z4ϮğdE��H� �	��e͊֗��!ɲ��xCL�x��I�����~w��+�~� �&�y�Ei���fi�צּD�&,:�#@�Ȑ����X%���������O��p�ƞ�m�[�J�,#�>���&8� `C� >h����h��\�����2���J��
u$a�ƫ�c4�<<u��c9�X�ؿ���r��,�~�=����.)��� L�茩XV%��
&�j|��} ��9�� �D��Q%㠁7����Z^�!{���x�Yc+Ͼ��4�Y�Ah��L�#0�����$��������iDgcr��t�A�H��\�_Z�M:������:�(�3&7�z8�`�����I����Q��۵]`��w͢9)iFV'�SH��]�&�Xw�Q���H�!=\��VrMiMe�ʠ?Ə$X��*�-I�g����S�L$�lo3J�>�-�7S&X�Dy4x�DM��n�U�ƼO23�� �B�tWr�U������U=*~�Cb;�1�9��$\N�H$�F�z1E��:�e�mX�u���g�m�<�y�|u���:/�~�Y���3�r���]Ʒ]�=Ν���R�Ze�e,�|p��sO�͢����L�(U��8:�(m3F��0�9�����O��Jc��K��1h=�k���̺6{�YyX¢��q��N�`�p
���4�0����3�+{p#��j2��E���� �-͕��U`"܆��	�@��X^9��duԺViS.4Z�"}����,�_LHkeW�r2��U_&�A��]}^�^N4���-�n_�Yx���'̯ �xX�$���{��e�dU��T^ �"F����P~�X�#M�pD5�!$��n�rL	U���{ӿ��3Y�q��|mks�������*����Rk�bצ�^������F�=ƕ΃֓��0s�*�>������V�	�.�L��7���������B����0�՚�S�-�2�!�zK�-6	fﱾRA�<��h�E6��pAt��w��v-� �Bv/3P1��^=�;�H������A� �Z�o�>zA�R�����$��)l��8w��k<n�n�#`�����@�.Zc���}x���Y�'_<��/�<�"�b����?�iމdP�q��N��S�B�iƀ!0}w�+�QrGk�ɻ$ۥ[���<#�q,�e#$���K��j�y
����!ĳVw�̛�K��M��9��8�O��+�X@�/�20>K~I�߭��6x1�¸c�_e��wI{�{�[m���uV����D&l ���5�����-5xM@�Ν�C�fT��|�ԭ�-�&��d�HM�;6�&~2������ԏ(TW[����~�֔���K�'z쬨sy����C�9�u	=��k�u�Ex����2 &��R֌�:���X�c� �,�a�O���}��w�x���Ռ��X���X�!M�hd~S�祫{x9lG�����n~낓oԌ�+��*	G�O 0����D�i��R1/�� �F}	��-�5d�� �H�d�mo[	X����-]o0�-)�h5e���G���w�?6�.�w�ƺ�DB� ���hv];\\��xA�w  �iGu�oq�|��Q�TJ�"��<���kG�5���ΦyY3�Aٜ�w�V�g� �����O'�ON����$|�,\pkpX�1���7��&��h����>{�F��q��s�5���a�@�z���~u�5V��k�"�E3���/�фt������y����엣� ��"{�{�f�c>�"���R�`�,yȣ��Tʻ���r]�J ϣ�a�ݴ� pA�8��7��U\}��9L�h�b�2�Rd5;R2�.���,��{=gD(.�"��Ƈӵ�W^ρ�{��5��(f�I��p<&��4k����7Š6$���U�|b��|�;�/��cOZ>��)֜6l(~}u�	z>�q�����X�1�[� ���%��e*��V���20��YW6��dw�ˢ*��V5GƘL�ba�fX�s�!�ʰ@#��Gj
�ZôPϦ\V��>��L�����U՞=mF��o�c�F����>:5mb�Pg�Z��Zf�7H|�fatW��^(�Ķ���qv�l�s��p�}Mى>X)�^4�sG�q=j�<MZz�x�8HbIE �f&m�6E[��z�f���\������=7TΓ,�� ����+5}~w��Z\�t��+�j�_�R��*_��9���^���"#)F��f�W-:�]�S��hh�c �6�N�
�аb��������4�En�y�89��^�|7�N� ��H���});֭s9>f�,}�R�P)�=���!*<����$ ik������w�l6\�P�<#PT	M�i\I������c��V��KB.}�;Ϡт���P����Pq_2y���qg��:�ncG��Z#c%^���� ��Y�-?�h︽F�-9����xju��\��a��4uD�m[b%��/�2Q��C������*��:�<�����>�)���]`Q5���X'�����Y��0�Ig7�ںJy�s_�5[���9yjT%\�P��7�)�&otM:���wX��e*TU�,?����@.И�)p��KQR����{(D�h�[/%�%�e6"f��B�5��4l�?7�Qr��^,��)uQ&O��&�2��uɎ�k����W����Hzѕ�?��Ĺ�y��Y�E-��*����U�M��]�� �#Tp����EG-�2۵�n��{�P �9�rK�Nס1*���u~��&��#D��!��	o�O�Qc?�m?�����	&���Z�lg}����Mt����?�Ӈ$��X�ԫg�N>�J�GH�?;X�<�<�0��hb(�^�;L 8���]���p��K��>9ZzB��_�<m�޶P�F�e�#B%�z���г��y2��+��/nzy,ڿ�p��>��&׾a������VW}&>%����f��Ԧa�Qr�b����gVз���#^���(m����+��y�L�qgFc`ß�Ra�J�
��?��Z�#<�UM�ùC��o��+3`��C�F�8��Eᵛ-n1bǸ�m�o_4䒱A��K��TY��!���
k!�?&�ݲ�E,��jb����Y��#@��Wd�m��]�}��a�'���u߫�z��G{��e0�`Y3b���jy)�[U��7 �t���ٿz��3ޱY�c;/��4�}�[���͑s��Uz�sN4����˷&��0�7�oc_�`���wj�E{���G�~D�i�����u�������������C�͢��jD2hE򊂍5�=l������PzWx/.��U8�[)
���8@�|��G�r,�U�u�	P�V�)�VVd�)�����goԴp�����ߡ��� �Ҡ�� �]{w

:�	ѭ��ы+`J�
�8��Z���5�^��t6�8cw4���a�DՒ�3�R�Z2��}�V՛ �D��qK���hʐ �W�Z��È.��4�����
#�&Å(�� ��䮭��?��י���<�C�:��x�+�߹�����,#�&�̫V2~)����=gKRh�)��C9'"g��;�q�[����L2���Ǎ�B�U���C��MR�Fyh��@�:��je,=�~6��V�T�ka�/c"���Y�w��!ս,<�|c{�yJ��[W�$6��f�6�S+\qPV�Y�X��M��	�J�����b��鉈��C��ϮY/�\�$X����i"ܬ{��*ʍ�Ñ�J�)�.�R��1Z��y���C�����s��H��b���]�����P�D* �(Dr�͏w���Y]�5u������><;���3�?�o����!LblA�##̓N��ʃr��T�yKF,6��.�D��1ٮ�[���恚��Q%48-�K'�%2��������^H^��]�̵�l�����٤^.����I%8Ɍ�]A�X�8�����x���wRr����=�_���D�Ds�z;C-]��>��ʗ���%F���>����2[�s������׿�J,o��J��
�����z��Np��2�{_�|�1�y��� N���,�7�BPj���&���@��Ҡ'�jc�jK�y��*�NA
�~Ttuw���ļM��\sS�ꮉ����wRx�K���h��&=�R��_龱�ԥ���-���,�{��R�rW�$~��]P-Sqh$� �h`Cy�ܛ�k|�/�S�~T���Q$�v9ٽP�
D�s�~��WT��TQ58߱� ti��g�"���0Ǵ��Q $j���c��̭����s�������/|�@,��.���u��ŷ�REM_'Jt�x��j���Y���C��p(?#v��F��l��{,beu嫖t�b��s�I���hŽ
H<ҔP�X����ô�b��>����/^QW�F{��#�����_��\���&�T`�٘D���*e$*O���U�g�1I�)�O?Q�ʾq�I�O]آ0�G�o�6Ս����Q��(_�yHF�լ\Ɉ)~��qи��nO�' -�:kxo�:߷b��E�t.1�㨧��¹�-��@c���Ϣ�p���&��X��x�e��o0�����#�������Q�����R�Z�Jk͗nDԃ�'���!�s�ک¸xe��+Lh�e}�y�]�pA�*�8�DAu&b�=`��,�$��׿�kx�?��i\��[�j ��g�c��	���q��O�\u9���v�#�҄��V�6��0��)z K�
j�`��c��-H����F��WW�n��T��S���:c�'&jl�rt�]�a�m�N��E;qܗɁgQ���dI 
�w�h1��@��<���
/�}��8���x4������R^�S_��}4����&�5�E��OƷw_��n{��'W����Y�ǽ��׎N*�闬	Dv�)�_r �ht��D�@����uX���t���^RW �����0߰}� ��R���!�)�'��2^�Ѐ�k�f.�##Y�/�Y�]o �w�{ǭ����(�+F���EHzx@��ς��O�SE!��s��̙2 ��̯��E).�C�ΐ��F���T��
n_2��DcI�FZ�ca�W�*�U~�~<ǈx#�٫U�"Ƶ����ǿ�d9{��a�#��3�Q�r��MM݁4��+�D�Q��%`�8�;T}J~�N�s�(�/��0�����FB$�M�~Q/���f�e�D���[�:7��;H���j����ZxYE��=�2��r0c`���?5'�y��_���rDo��X%��#P����V��_Q`���N��پ#q(�Z��$ �)���u���&}�����O,�l7Q�6Yc�i���.�Tc�eo(�p���Р�xW^��k�mRQ�K��0�6������Ta@ϥ����M��%�8vJ
�?��Z
h�w"�=��63v�|�k�s}�=����������$����*�j���(%d���H[�J;��9�x�k�|�W^�x���d��nUYJޜ�����%!�P�L����U�W%o/$r&.fId�{y�V�7)X����0�G[�����>	@�q:���O0�Ŕd�r0ꏽ��{���u'F�#����ù�+��oi	l�Cc9b���j�T���h	#��������l|x󘳃9���æ=�m�0�b��d I��z�ݏ1�U�E�rbD�;�枺����(�-�ҳ����:ߩ]0ňw�4�e�>a��Z%tR�(�iIOf�"���>���~��O�D�P�d2�)��7٢��L ��y�['�kk����X��,�x�3�i�c�=����$)!4��� @�w��OO�%2}M���i	�va
��?���Jp�J&1Î|�w߾U��J�Fdpl" �l����6�M4��(�;SN����;��9aBɍo�~O�6K-���,����?�S��t�ZN������1d���>�@��r\�^��MB�`�A.v�I�V	����TR�fʝ]?D=���Z��b��p����e�c�B�p�H���m�
����g�7_���O�3ª�{&�i�%�c��VE�n��Y�W��1�*.*CHk �x���b	j��T��X��q��8G�p�&p��op����|�T���v����C&*e�a�75�H:���y!� ���295KA����$H����E�یkb�-�ծ��u�����l�b��5eIVw�>uQ&�y�&{�����6�8Ì��uL=|�*�B t�뫌�S���
]����8��`⃩μJ�z����Ê/rH�+;S��'�X~��%����/��4��"�
F��#u�����q�����sb5�ɩ?�ŔژY݅�&Jiu]#2�5 W}��c}-�jR;5��B���j�1��(v;���e�S�;P�!��� �9�2n�^��YP�?��ȹ�@U"�P|5~��� w�M.T��.x�A��Ğ�/+^�y��,E���0^2=B{l�X�v���r��a��5��&Fn����v���Qت�t���XͿ���Ϸ8U]P�l��a�
b� ��-
�u�hWC�@����E�%�L�6-_�8[5ѕ�_6 �6�D%F$������0ȱ#F���Yc�!~ڿ�T���ńo Y�4�;ӎ����j	��y4p
�"��+t��HrRfũ�G��{L&j�PsO��̴��Kѣ�4��(^u���)��.7v�: ��O��8�f�}7?	7�����c���z�FYi q�/E�<���P'�6�ƾ�/�)s���f>!X�ͺI�<�&A�&p.�3��qސ����}����l��� g�ef�`�=)�z�S����We!�)�e5)C�ż�q��#w��SO����g�6"7�6i�5�!�3���~�-BIze����G�}��x�UJ�M�;�M�9��6��
FS�z5h�I��.�)�{�د^hv���$gul��*2����Y�� k�e_2��v*��Z�C�����*k�m6q��Lu~��1bw��<���������?�|����*�uK��h'Q�4^�� o���b��U(Q��,�y���8��9^��D�`Bċ��&t����Ӿpt0I��Lf�I�=�*�(+UBI��ѸRR����2�&*�,���~�2I!�a�@�ÜeP5�@�ķ^?m�-������ƹy-h�o�͐��+/ѧ�ш��E��ҧ�I���*q�+�rfWM	ld�f�lkL�"�*�Z~9sCP\�	����Ǽ�I��o���dVH�3i�}=���ɤY>�`�y�[9�!�;K�������˥Hć�Ԥ" i1��䪺���kV_y,9����ߊO�d
��=_�"XFId?�9�^�e9Ƚ�.���bܽlQ,�.����T��T��>/�͒�ڱ�)xWٛ
�k� 9Y���;��%����U���ʭ��dM�D�/�㎠*l(N.cj\���� 9�m#
� ����j�P��+!� � ��]�R�L��	7����E,�����Q���!1�n<w#�$��]�\�S"xV�a���_�f&�����o1+P�b3����[��ۗ��#J�!�jS|��ҩ"�=�a�w^c�6�31>��q�9����p�6���XE2��"��ۋE;)1�7�ɽ�N���K%�@|ԧ/�K4Y&���z�f�So��Ed�)�Qj���%���W�m���ig3�t�a� �7Ke�M���VlG-1�k9KM��L�3�x�Cu�$�!��<쾏J{�����ySMBPU�l�b�����ǂ!�#4�A�37���(����:Jj�c���db�Ôil8�	\�����2]M�3��>K-B-�9�Z�3����|\�����?���t����pM����'�ї������}:\A�p��ߠ���ϙ����!�9q�vL���Ð���&ɮ�So�1��M��л)Bk�ll7x�W�W�bCӊtT�W����{V�Y�鮝����<�!S�i?e�3�K#s^�i�y��;����%Hh���Ŭ@=+��{M�>��h��on"m�(��� ��[)�B�[#F�H�c�W�֯� M7��V4��ع*"��v�fv����V1����Śfbfk8���X��Ҧ���?�}W1��\���y��bqh�1LtK��+�"a�lޛU��t~%���t�T��<,֑�w	c�T���=%l����<�ڿG���e%w٭�v=8&طY�lL5{���C�0�:	�땿z��hӥ�\c/�#����2���A��~���;F�0�?�V���Đ�/��.�%�noi{�~�K�J'�Ze�/1��Z"dz"�yy3�����f�P���[���-1�m��C�k�"5o&ñ�zcg�!0�����e�˟�c�f���Ƞ()�����=1��D:��!�6w���91y+F��E�\�3�㨞�J(��T�W{)�e�k�{
��ʈ�=Q��A�����>, �, E���T0}��]�zc�s�'3� U|j��@�F���y%Ϋ�z���(l3�/������ a'�f�KK��a�C}S�,�#���Y<�K�'����SظY�����kg��Q2,�rU�x��+�o�u��l~#q|3ր�YT�#��U���[���DU���.��G˾b�ۓ/���{�'E�]�i�i"��9��-���{O��,Dg�n����R�sA*B3�A2�4��|���A6=U�@�"��.��n�ǰGy���kD<N�9�`1��w�J�B�.�(�e=tm_��z����^ܢ�ܯ�ϚX��P���gS��"l�wa��\$�I�`VV�����i08� �j��X��6���h��K�i�����8�p�p�N���'t�v�sK�
���۰N�u�3�*�1pR��1]��������VS�2��v�9*�]���
e����W����4N�'�2"m�M��M�zk���>֝�H�� �Ԭ��Q]S>�a��ȅ);毑����Z[Ց@����hȮ>o<�*CK��}=��x\w<�m�Ě��2}�xx�V�{Eg�mQť�2�O{6@���x2�-�u������V[ˈ+��aR����4x�H.��>2,�A9Q�j�w�˟��Og�4�6���o���޳����73�f������Hw�s�ϗH*X��FpLn=��`��������D��H Ȼ&��`{g�$B�:�~�a#sʑ/��&,>c���� JC
��GoF.J���kf3��J|�2�+]��)�h\f�=��4�������:����Օ�e9�ڟ��eHԲ�y'6�&���Re�B�K�,\ӴE���~��N�n�Q�=&�>��e�N�K?ab%9���E�'~D,4$�j�����s�Yw���LL�V�2%��&�BɠSPA�GLz���(��G����T������$���=O��YEp�-�ʜ/f�(���O|j'�~j��jc�xп��ؕsU�۷����O��U4�8i��;vu���I�O��	)��0t��C�:��?�xs,�]C�#]�*KP)��-�&ڪ�����9��)����b5������^.� o��C��H�/V�Z�� ��7p u~�udv�K�Vj�isr���R� ��c���ۼ �y������$+�Vl��q����K.� �,Sn7�7�F�g�)-�EY�wE�j��<4��'o��<��)�fZ6E�V�Q>��ppA�fC�ưo޻�n�J�,AD��&l-ES��x�������T��;ѩO�(�1~����#��^;x�����[�v�L�-G
v����ta�Lx��	�� ��ּ��lQx��(������ƣ�E!�~9���!|,����A�����Ӂu�̹�s1��� ��B����[	�٫��4�xbӝ��')WE��Q%ĕQ���Xh��cx�椫Nğ��7G֠��{���5���#f8s�ƃW��0B2�[w%aI�|��
�9�^��Ϩ�y�p����&Ƿ���`;��S�?�Ԯ&"�.S!툽-���k9��FL`c~���zW��J��9���.�*�Å|��&��aJ��Bu�X����էq՚���g���. _�t��T9�U'F�9���S� *��=�_�_ӎw�W���#c;N��&���uz� �/���9�Jn������ƫ4��;�?�=���Dk?��Ie�����+
h8�,(�[���bh͊9��� ��s������'��˿�͟�=3�u���[���$�ߊWd��^�,���DV:������ln$�=� ��8�� 7-G�@�FS%͏ꓱ5�!gTh�w�ė�ڳ� ,�,>�4�&U<�)0�#�=���g�:����{P�o�6�b�=�Υ?��� B���*��T�b���1�l��{�3Nx2�;q��L�[
y�{����n� Q3}|�tߗ��<?�v�B�}�׍�x�R1Њ?��3r-�s�@�+P���uB9�&
Q��읏�A����$��X�Zo�q�Եұ(�+�}ʺJ���Õ?`p�w�4�-���C� ����\�c[�;12���IM��AK��; �q�Wa� A��w|��3߅��:t�]>��ܞO�H�N�B�V�U��K/�B�1�nw���{	��Qǉ"��q�И�\B��5�,α� I� a���[�Ml�I�צ�N��{��=纺K��"3N߾o����^HAW��OY7��gDP�=��0OF9���n��ʫ$�=3N�^׿�c=��oe����ٵ(ؓI$�p�Gj����X�Nr21r�l�b8�*�_P�7Ҫ�c��J��ɷ��&r�ra�%
�tE%i�s�$��[4� �m4*v�Y;F���8/���̼t�#�D����-�l=Pv�$�[#��u��2j�l�k#�	�>��86����-�e�0K�Z�$d��MwB�`Ad����j���Ut���PB�F����z{f<<�L�w!Ʌ�Ƙz��3k�vc��"����*��[	��-�R	�}��4���U���v�q�3������i'!���[E����R}���2���c��3l�Wm��xs%��ˡ#�ʸՑ0�Ԟ�Y�w�s+���g��u�"%�
��l�B���'V)�C%�P�~�q��Y��>��+$�w�z�!<�ַ`Π�5,�\�)�V�z��.n������B]��׭�G�ߞǞ"?�����np*k�S�tg
����O}��T�@�!�IF�%y��K/Q��;V�4��`<+x�r>v��l�,J��6�6�>2Y"��c�TF-����oR�L(�҂M�,�	�p���R�����)����:o�;����`�}^���A*�&�Al 9[�TL:�Gٗ��.��2*����*"�L&�[��sC@�<���J����/��J�4�آ�Ox������ H�~5^k�5n�8��3��[?���}�ܫ9VI�}���\��(�B|�|�iڒ�f���L&�e��������� �����S�h��%xd֥��q;��YeA�O��q�1`:��q94��nN�s|EXd���R �ZP�S�a�޷�w�_�*8�	�Y��˅;T�U����fw��aQ�
5�S���� ;l_�m`���BE鉾����/Y�����j4;����)��Y�8pjh+�����0�}�EY�Z�n#����MwJ�/=��}�C��J�is�ǬC�/���'8{V^��>�NՖ�(r�1f&��m&��mFW�A�.bU�3��OI�L�Z(30�G�;<�[��Py[��[�����K��I.~+����|L�G��j�@q�����\+`	�[X����H��l�whM�f������?C�8��C������7|���i#�0�����0��閿K�!�:Q2������:�Q��7�8����E�1^�IѲ�%�?�^ΡQ�C�k���*n:����T-P����w����@D�����;��5�w��2Ӡ?�(�ʐI��.��'�6)� �x('d�(J4�D�閎F�b�l6]���{
�p��,�u�1#�H492��`��P�4�NJ��{.���FD��5��$&mХ�Gvy�/�ޫ�J��ZФ	���ݹ`3d0 /7�X�VS��0ҝ � ��ɻ���{ah]-6�G��/H��������0�F*�o�U���W�q��_Of�qy9���g��ʝ	YO�!�\��
&ǡ_�`tf����<.��e�e�U��9�H�{#H3wI9�g���"`�8w�G@�bG��5M�:���|z]�L/�\?�G�GǺ����{�=�+Y��;�Gy{�$/:WO��bs�W�?]�T����`�4��z�"� q��n�C�>9�P�6��u�_�:��B?v����)�D�ebe�D��-[+ubM6}�Vͤi�>O�+ۅ1㩮��iH�Jӷ��:�1Qn�"�lc���/�\�tCN�C]mW<S������0�E��
�m)��Zt���3�)�a�M���g���4�%�d�(��;�4��A� ��J<g�a[��˻����+Y@ꖚ����3��� �Ǎ��B1	_"rK\=�:�?<��t)2��*4��X4� á�qϥ.��X���o�
#��rV/��]X`b��zp��v���|�xV�����,�T�������<���s\�?e�Qz��3�a�́˔͚�@!�S�̮�A� /�x�)[B��x��aXwXL��9��t�C���%-�~Z����&p�PP�u�a��5k�7ĘQ��D���m%�Y�X�'��V��Շ�^Z+��^oI����b�
I���f���H�r��lO� &������}�k��fm�E[^Yo�5��"T��2�;���>�2�F-M�f�N׆��zG���nfbR��.L)o�5�����k1�[+�9i�P%�A�訑��E ����q�K�+�+�r���)-�$�z��|T�GM	-��zFۇ�ςVJU^'jw�[i�ҏr�[]>��I�0�"�C����im���C֊d��b���I{�l{�UN�Q�6���/Oz��{��]S�]V�����;3�<+��l%[�gċ��|𣊽��K�!Ăd=�eXf	Ѹ�����B��H��x�/��Xb��7���u�q*�x���c��Y;�_?�ȕ���(>b�#�'��&�r�NP���=/5�m��"��B���c�Ù���X�Ƈ�u��䜡k�4��sux�@��G��#�����fЊ��)�֦e`��������f���
��e�_���a~��{{��ԯ+�[���_t�/<�Ge}/&
�3�C�᳤��#�8g� �^N�;p��X]���Ѻ/*2|x=��?�� BI����j=�1�ň�&�*��O�߫L�c�k�(�DqJW�v�i��+�-��m㉜|��}CB���7_�H��X�C�ho�6��-
�P0���!S�
AJ��a�r��,z�i.Aå<t;�8��&�UJL��w+^��a�R��*�j�ǧh��!��eo�㰣�k��nP	�Q"���X��(��W�~�֎W����X�W GL�qz�ͱ8%�t>��)0$A$�����'hx�W���x��-��A�l���_�8*+ſYێ��\[��B�w��t�V��ck։��`KL2Lz�[��Ϋ��bk*��^��}W�(�i;3��u������0x{4���s��M4?��A�+7L9D�Mu��u��F��l��"�ίC)�������Z_�0s������v[#v�,��n�P���?�S�zv@t��U���^�՛�+09�~��:���MP�}'�K���h�b�SҒE<i��K���"慛Q,d�ԁ���T�����s8.�匫�b���Q�4�Z����x����hQ�r�P���Nt{��P�yY�ϫ�&m�����c3[c���P��r�����Ax�(�./��,�$k�K��h�e7v�R�N�6�-|�,����2��~Ȃ'Q�b��7w�T���Ӽh���"�@ .�<pA��UƼ�XLOG��+���Ҍ
6�A�Z]�y�&4qKp ~��^�̹>�^��`Vޝp]]F�0��v��::�H��|nF�n>�����El�1_�����ڦn7(m��_�dV	F�=��C��;��������u�[�3�,��e��8,+�A����X�|���ᜫ麏sƩ�
M�3)VV�G�[��K���s���x(���Z|��w�Bo�?�`�)�*R��̺x�6�H�����7<@ږ�פ��I�f�$�^ت�(D�3W��Ep�A���D��ZW�#�	�lǧ�`�	k5�k��6��F���}�� o�$�"nJ�N�in,��㑿O��3Qn�����D&�|����I{�XPZkP2C�s�J~��i�H��ӯ���~2=�发�׋%w��`�G\yuh[���U������Lo����0�6S��!+yclQ�ٲ{��� �ޞ�5���04�R*���"���s�1�vUa{��T��rz�ำF�����������F�0i8�[����!�A@~�\|Be���׷B�lgĪ���U�a�y&��$����Q�����(P�&4"���e�Oe��ɤ���'��3x�Ai ^�	�U�2��7.L�(=e����?����E!;�����}I\�8�ȯ>�_���*Z_q8���|��(�!��K�����Ǥ���YN�u�2/Іv�7)&�����nβ�n�z��K�TЃ��̀Juu[O�@�9 ҫ�%;��D���s�I����;�%������;��Bu7�s�ă��*����*iKOa�{�T���@�)�8Xk�E�F�1�%Y�b(Nu��3�c���V������ ��.�J~�W,�`��#�h��6�"+������(�� �G�-������\I�$5�6)�]������MA�Ǚh�Jb���9�R[�����X;�K��\�J�_)��0pg9��L~U��(�/d�s�,
up������-$d��%!qrˊ�8Ka�tA��h0���&���̐�b�+���R�x���a��L=?bDdr�,W<W��i�����s�[�9B��b�u*X�F'b��נr+i^Nk�)�Q26N?5�m1� T p�ȣ���>�cNo�ޕ��b��?v�C�+0.V����I�i�n\��5\��譻xl2�(�xEY���F�U��!"32�)x��AkGp�e��O(*؀}��-M��`�I�<"!�L��mq�.y��%��&���c�`|%�$�����ZC���{�]V)�w] ��^<�����<y
9�@����0��y$CM���O�%���HL�H_s�^��J�o(w��\��_Z��},�Ԍ��/;�
�/�9��\0�5x�Q5�齭j�3���*��"}�ܤ8�/7�l�͂a?A��6b�L����~X�?���`g�@'M�Z�yG�����X��w+��}�+v�V�WՀ�����λ��tc�׫�%Ŝ�PT���;����P'�K)ET��f�`N���֐3XK2}��Τ?"$P��"G�:L��n�(�^2�,_��M�}�;:y��
�P �U�;��ˎ@�K��8��������gͥ�Wx6�@�a��efǎ�[�+�<�@�h`�2v�� 7�?��������4����@w<�Z��Ym�t�����$�U��Y��9�zbM>�@T�,��x��d�;�|^��S��\; �r�ı&c	�tF��=�\ӷ����m."N���qFVA�(��4�񝦂^jY�P6r���ǃ�s�@�xV6�|=!������q�`|3#���Վ�l�݂*�Y�����;�Y+��B)���bxK�r���1�/I�}��̵AQ��\�b�ܐ���{U:���OzJ����c[;ra#;�aO1( M-�.�
v/)�6�ʟ�?��(��spS�G�Π�ܓ�8� Ӹܲ��	�A��*\�� E>���`'F%��u���%f���������߄�*۱1�6��Aӟw�q�+�St8��)Dj�-��S]��;���fO�]K�Qd�ud���i�`:>R/{�a�Zś4�b0K]>�u�GSM5Q���[qǤkmN�a�!�v����קE��v�h(>�̝q�-a���g�3��^�}�O�&�V/������]�*�؅��*#ģFD�{�)���r��n�xЯ���h�Xt�b�Nr��L��F�P��iSK+V�N��c�4P�;�64Sҵos�E�wF�h84)���O�Z�jL)�k�XB� ��Sۭ�׊tY".�ph<� �Q/���
N̨�B+C�X�Pz�Vx(���p:j: 6&@&
nX���:�]���������f�/��Ȟ������H��?�B�f�(�Ϟ`��)a?z�+�[�/����_��G9z 込�{�D�וD�,R���ŕ3�J;�?j���Gg:^Ð&4��ml|�8�V���:�N{ӊ¿��if)k�E%0�Qv�O*����ߩV�ҽ��F)�Y�C����L��=� ��G�$�4bR8��$�a�ʣa�:e���BG�6�rٸ��	��>�l�o|�p��m��TBd��:�&�)Չ$�4��l���clcj<�((2�	[�m�d?�d #�"8=����wyCapt�[�什�8Z5��Ԋ:��#�6C
�������|ԗ+Y� ǧ�SR�5�1P���Zn�u����r�`��*��܊����Y��I��{�!��z��q������CU�!'dJ��`�z�7 ��`7/Z�Q�����%��W��m*$֍�
�c%��r��[y��*�{�(�!E���*E�g����X�CB��f�s?��V�jNv�[������^��4��-HC���놎*r{�1�T�p�WO��g�F�5���y'�KOb$�B�qf��a
�b���7t��C���9���.gO�� ��iW�/����HX2y���$9��B�Up�����K9U�Q�a����,4U
=��Y4�# w���jƏl��8ԋ�ʰ��eUp��=k�&�v/V^�H�W>��{<�Aޙs���aزe	��!�?f��p�+י`��Ѣ��_-�Y�1�j�yݔ�Y��rP�6.�O<��yi/>f�W������<"�1�� �ߜ[�<u��y�$gN�)g���C�3z��O�3�\�N��O��lo@O�_����[m�dYJ�9���k��}����z�0�1/�C7
_�P���13��W�w�3O�d�:e~W�*��J$��o�[Y�7�j+�?&�뾮F��k�+n�H(�K�WN�0ׅ�k�R.d�Y���ൡ�P�E�.�u��B^),�B���^M�
V������h��b�k}lh1�S�bfɁ�=7�wo�	�A������1���cv��d�IV.��5��Ѵ�_6��/+}�m锤��W.�_��^֩��-��E�Mw)$�)�ɬ!����9�Ł�_�ڟ�2<&�1 ъR��&?U�(�����y��P*��sN�Ø��T��I�I�A^i���}1�ZY��x8t�n��Y���k�Ƀ����u������������SǍ�0(Aab�'�_a6(���!���WI���H������ ;  #{��h�+-jH��6@gA�I�=z�D;����'���` R��,�)�����C���*��Ɯ����,$ �mV�ӒQNАF�$��V�B/oU�D�V���8� �[��E*E&_NiЛ��N�eW0	�W���|pj
��`Ӝ�8�ԗ��FT��t��K���̐'���vl/jV�#�0>X����'�*3��k�Y�$�ȁ�0Ų�\�tX�A�^u������4~9�*���D9�37|KB���ɾ�C5���չ��΁pS�r�༴9�ڽ$�ԅ��Uҙ��c�L09��^�*�v܍� ����\zT�5�ŕ/�R'�A"�yj�MD��M&V|y�# ۋ/�ӎ�%5��S�Ѝ T�];hA8u���B!�9	��߾�D�qK��^o_v�[� �]�a�ᵈ��z{o�Gn(=��`���)�7�� UZ⍘\�X6:��Qy�}�H��BɆ2��(�/�~:;���v6��{����:|�3БNf�sX*��4<������I�|��d��X{���f;�ǣý��hH�s�'��f�~�u�O�K�m�q�)���3a��j��8�� 8ehNv�x��|F����*'�,���i^��sK��b���%L�Υ	UACFWYq�g09By3>\gQp�k/�
��+$#,}+�Sb���0�J��=i<<"k�l����؟��Jeb�������K�o���̽�	d��nc0B8�D�ES�_�R�(!&ͺ�nX�sD��z9��ܸ)�������m-E�
�뷢��p��߈h��.�$�}Hu^msW&�6_��L�� ����;�4e77��$�f*vҞ��v2�R����⤴j�i��f:�@&:q'�'�CY�������@%B��zk0���-�s�v�!pK5�zq!��[A���X�!vb}<�{7E]ߋ4兗8ݽ���Oغ��gW6��U���3�@^�����!�%�6�x���Wӂ�K�so�F�A�y���Ͱ�j2* �m�!B��yz3�t���>E
�J�?�=�~glS��u��������T��d.�#���94�ns�˜Ǐ�,mo<=
Ogo��n\�忨fZ�$���Z"�7�ϊ�Z҉���=��Գ��rY��;�W+�gT��k䌳;R�{��x�ʀ�U��	t�_�Eg�^�i֜<���o,��|��g�:��^�p�t��\.��:e�i.��z�ʡx�ڃı�H�b��� ��~ղ0����~*����� Eg_���8�#��=!X1R�m��f�mo��E�j w����>6Æ(B9�kO5�}�$�@q����w��>%=)�^i7�> �O�	�T��(���hjL�YF���v{�56?$�iR��#��IQ���i��#X�9.��,���O9���K�t1�����:��HY??7L���`ݟ�AV�D[V|`�ּ��]�V2i�E���y�g��rᾩ�J0�Eҟd�\��P$Ҏ���:����c�8�ˠ�-���]��<D����q�ao�L��L��õzAJ�N_֤e�qٿ؋+Q���ӻ�3��	]����J�%�821��Ǵx�%[�� 5�2�65�"1 2.Z�l�j)r�W�69��1�Q
0V����(��Lڊ���־X�".'����g��%�3��S�Y5f4^�B'��S��zM2�Z�������>���8�oϐ��ҕV�� �je<���<7��<.��9���/�oF����F�,�M���s"\�̜���D�v ���ȏ�H�����5yFa΄h���������@�ÎaQ/eq?{�5�+3�-�������)�XA])��9o�/��I�W�I��lE��^�.�9ܛ�`�sM]�N.I��4O����Kj(��+.$�#��/�^lֳ��-h�S8:k�%Y���2#"À�/<�(���#��ao�{�s�nj&��5?)ǲ��Gػ���į¼���س�ߙ}��i��keW�I-�E3��9L0��2(���+jUQ�-g[s)P"�HҬ��ߑ�Ն.~���_�@F̥za4��fz*xllU_��Zm��3�K���Z{�U��dF��F߁�2�����xj�d4��?�h�T���;@�?��,�d0P0"�~�~;|_�C��
\��(0gb˰Yf�s�LN�����n�q�l��� ����;D8�O�h��"���8��Z<��)��<����{.�pI�i
:��W�u	$<��||����NF��N�}X�&��e�A=;q���3�i���U8v���3�u���i�I����T�S2�U�?���-�w�ܔ�'l���_u� �]͛ۅφ	ÆD�����F�Z��(\j��x���v Q\7�G� �h����$G�8b��)X��"n�z�hb�`5��e�T�V���P�6{�怿��m���#k���l���x��j�%Q���t����B���ƿܠ���b���ku/�h�)�<MMFu��GꙨ�yF�jE���@�-,��2���m�Y�� {d��t��.°p�#M�6�a��2#/�[&H��B��e�!K�������	����+��A�����w��� � �4��êc���!���C�ĩ�r�~h��Sf�1��7g���%��%ĵi�bou���� c\\3�;K�?��	�?�y��ɷ�=�if�,/*E����)*X���͖�r� D*�}����.P1�5S]����O~�ݸWD$�0u�y�P5��@��w�ck��َ�/N�f�܂������=K���Q�~ ��-�����qJ�'�4�5���
J+\Ɍ��;��D�������O)GБ��#,�@{����M����@_���g8(�@�"��G�O�E����l|�hoܭ���*�����?��B1[V����rg���֑�/��H�9S�B���60'zB�:,�V�<f��q�����g�-�`��@������؀�9�)�NE+��a=V �2�9}����`r�um�����z/�C@8��Љ��h}��8��)1��5��8�����P:��?��ZPn�Tq�߱0�-BPM<�p@�v'�I�A����T؝�%�P�N���C�# SWU���{|�������n˱{�>���u��W�l��555�x-(�t5�����<+`�yY����H��WE�Y��Ke?�#����s��"<8�4�6ۈ�����gOm�ʍ1y���bbJ��^��1˴�+k\������+ �SK�X}���Pk�K������7���'MP2����l'���p-��|���aA&t	�Ĥ���3�c����7y�9�jj����P�F�o`�E��V�j�b���9�.D��� �R2ǚ(h�(�LQ͒�f��5�O�Z����Q���_��|ώM�A�$%2LoS�R7��S��ڎ�/)�ym��#���Ǻk(����m�ׅ���ئ^�� 1�<"�i>&riK~GG	3\��Ԩ�Zp߳[o��n��1�>�����R��&��]rjj@%,D�Vu*�Fg'�6Բ���l=������?�Cf�W�����,D�y�O���&Q�L��m}g� l���P����1�Nu�n)t=ze�Ύ�&|�����R^3�ib"=��X����G����%��;Y/�p��1P�:_
zë�wt�G�
̑�j������|3p��<�8ؘ�}{L.����&�nT�V-mzj��O��)F��?��9˛*�Ikc=W��S���a%��)��Z�Z�;c�0��4vOJpt�����2�	;/jL4�c�R� ��)H��c���Y������za�ǝVkZ���J~�'.�T�lgC� E# Q�+3}|�x�NHT��b!ş@� ;��YW�JҾ�Y��j*���8y�XAS�.�P ����Y��j
�b��i}���~����K��	�qn���{s���՞h(tCH.�g����A�˰ͥ������c7��^v/�
L�/�"���^��$���i��5h<p�� ��:;2 ��i��ˇ�H*K������=��ǭw>�+��_��?�+חVp��%X�J��V6�c1�b!���eq�D�m��&.1tVo�.�\#����Z3���2�~�s���6���FUu U,+F�ī�u��M���!,�GO׷������0^3Lv�-*d�����]�S���V(�����->j�2	���_�8��vD�)��!�V,H��O��������&r	�Y�aK��M��jT�E)� �E��a���j����ZR����yh鱂��6�e�8!S�Vշ>T~	_�h��5:s��.<hIk>�r�{c�ZBӢ�4�����)��I&E���:��5-��痺�ϔpN�Ť��I�)�m�n�XfLp��~k�p�c�H]T�Xc�M�i���Ё�L�C��go[x�Qo5��������r؛�ͅ��(�D��7�T�#�EnA�9����y��p1�����! �J���cM$F��B�p���O�e�o���.�"(V�Ip�`MW�J�A�-�5�����OF�|z���g�Q�ғ|�Ge�����v�I��/�AT�fHZ��j�g�s$��N[lM�C�e�U'p^�Ah���2��	DT�6��b���aWS�@*��ߖR�t��b�w�,��$(G��K��������D�W�3�g����	1���n7�P�["~�)�R���?r�����!��ԗAK�s$�ؽA����-��ţ�ܖ�&�99|��l�ovЕ<�ݢ�,���3��X�����Qs�5a��ʠ��U�sB)J�ѱ���������&�A;.�S9_��:j����o�\QT�<�<��N5f���)�T

i���2�No�)����
L�O����2l���;i~w�-���sX��;蛟ݗ����+�U�-d9���]vמ(�<�hK�n��8�V>FC�Pѭ1@���G���!;�&0hg��c���H�^9$���&�)�6� A0����=	�_���'b��3�}��e�Z���h���������WM��-�d
^��p\��[������fO�d��z��rM�w���v@Mm���ОG*X�M'ֽ��؞�7ҝ��a�IJjg�:ێk5��^�]eR�*x;��^��R��h�A���(s���"���8_u=�����=t;�#��_�5}���@�.&�������+h���;���t�V�T5�<�����hg�S�1l�%F��������Zi�����AJN�|Iؖ-*If��@��\b/�Im�^]sG-&�14�`/�W�F�+'����T�x�倜��ǣ:�) �,�9_hyW1�F
��~�Q���.�f�Ƥ[2�4c� ͐�V��^�}o�L]�j F��@��H��d�w����U���Cf�`(����0w�2l?4�+9w��pg�Њ���Z�H��u�(��b�$6���+�F�(ӵ���)�Ul�x�M=��2Ν֬u��K���T�6o����n�ճ}r�/iFaH�����W>T��J�Dh;V$�Y!bs�/�(�\�ܫ���i87��nA�;�B�,z�˪zh��?�Wj/(��>��LM�rM�@F���(c�d��Bi�/�qRۻo\_�Htj�x�D�nq�q� �_��Ho�~£2Å�bb-TwP|�}��/A�'\��^�(�����ϩ������9�P�A�$颈/m��u:E���~0	's+���L��i��H:>���:;�G��_(��Ӳe�w�L-8.�$�9�4�sn8����r����P9L��w	����+�K �Ԓ�ۛ6�{�@���Oy��>�m���<U�},�^�/��!q2�
ې\����`7�� Z��Y����)BK��JS)mx�4�������5N�O���;
U��Юg�Q��4$<���I�a������Rn>��
 i/r���_���/X��I^�vT�[���+�z��r��ʦqp�/���ҩpl�����%�c�+ː�b��N�j���5eM�$�)���sZō����˩!���1֢W�+�a�e�\���pá���OB#�ySɈ�mY���J�V��]��Do�F�6�?�S,��A���U����Lr^�ǿ>�l��e�vR�fv�)��
\⢴��n'�%����f�=~ ��������YO� �2(X���� �	)͐s��M��@����8h
�Քp��2�I��7�,�U7ߠ,�l��3C�?�5!k#Rf��jW�{К�;Uߙ_�![׾톟@�B%�a}�D�G��U����
Ҷ~��l���V7�=O�$Gݸ�K_U�G_f��3���eW(��XG+އu�0�9y��A�ӱW*'M�Ҷ]���zֽ�^� ��"~��Ԍ!ُ�g�_�wi� ��eF�(\���D�n};���&��Q�d�����(���r�1.���9^ˑb~���+	�Df�	�?���A䲷�� ��}I�yfQ��ĳ�ў���NM""������q�hu�N�_�������g��P)3~tC'C,x��w���X{h�N3������	���(���ҫ#����4vY��-t��w�Y��a�\d�ŀvd>��Y�݂)��7���k><��W��{3֠� �_�g���?�U�!�8�8����=��Uc�MF�d��.�s㺍s�DH�%\l���c$�� [��1�(ԍo��/-��zQؖ_/3�`��9�ɫs���J���K�el8O�pGn�ۯ�i4"ype��]�M�}1*�HѷDe9��m*ہ�N���²�[�a��^�K��p�L��m���ۀ�h��-��&�2�v{��f��Տ���q{��2��Y�4.���Tf����;�miO���r�gӰ&4B���͟��>䫃��d�^�$a&�A���
�A�з��v��тb�g�P������S��\gRjf��fd���	�2���"#���R@��*�eZ�C�A	�HE)zM~5)�ER� N}���5�K��mam������j#�m^�k��G��]Ȋϐ���f����/X���e��N��DP[ƕ��,M��oZx �]3�-�xC�(3yԗ��������d�5o���s�&l������׷���c��C���t$�AnV����:��D�S@g�14��ǂB��|���oQ�b��:B���C�/{r�@d���(5��}nj�S�O��3F����e�p��#&ޝ�C��2e� ���ٽM-�*߮��I�m3��RK�}X�HM\ �ݜm�U ȉ�A͂D>�����*���x�v�٨3�����1?�K/m�l}}�o�@��d�Mß2����mťd��r�ul����w���e��s�X�h��`������և�T|�{pkV�����H���l�1�	�f0(3qq}��X\���6{�]�4Iy���<�[)9��+Oȃ�������(xpa���57��{fe�*������̮_/���P��XaS�t7,B�'�Y��������Iޟ�aU�e`e��Dp#���\�mNx4����K�R��c��������h�u�a9� �1�	\<֨�O�����+c��d��܊f� �*��~��0������l��[~�3r��Ҡc��1!P5s��G6�H�!���w����Ơ/~��l��f����?�ͱ��a��&�e���&:>t��<JOx`�X�7Lk�^0-��?�wIo�.�b§�`���j��^I3c��eQ�"?�0���ˡ�,Om?�fO&.P+n&��N�,e7�q�_!^�[���H��Cu�^c~�q�Ӥ�RRFHsx+���i�!oxoai��v\j�?Y��v��#���O��؇���`�r/�n�w�iߟ�����q�eW�^�����J,���WO)|�-�ɺ].��$;	�}8i�հyY21�L��dbHZ�6��j��v&E��!$��ړ�>��R�I��N�������aB���e�C�m0�!�1&@�bK������Z|��b=��Ӎ�؋��X�y q6��.{Epa���f;�OD��/�n�߾��P#����i�ؖV����ٗ��n���+�W�$̙K����M�p����p��a�TD<��D����)�	���]�F���S�[���c�R:�<잢�m��دs}�|6d�_M��-P������/�p
G�Ilg�%�"t��ZLd����+�gpc�����;���%�O��M��=�������f�`v�#��!�T���F�5�:�*{�U�y�=-f� ����rq&I�B�+�S��(�{��@���Őˈ�#J�'��|��g�1�0L-	���?���	���5)��������SRl���_��2� �R{���D��։�V��\m�P��(1��z�m��D�YW2�|`(�v�f��5�%g���������(Dt�M��5)ip��{���	+[��f\�о���̨�-�Y��~�5�a-[�uC�rӖư�z�_�]�v��WBľ�W�ł��d>yO�\�k���[��/_<b���i��lKFV��z���D������
<��q[�
H(
�5O2���ˡLO����L�F�k.ᳮrz{Y���T�4�>�Σkc����5膾��Ʃ�E�-I�IH;�����`F������`vJ�{��])�����B�$��v8�CS��/��b�4�h�\v��X_]����� �O��{���{��8i$����%�oM������/�w��y�͕�^��-'8>$��:���KK�.����$/���j��e%l3�H��'^c�X��]D��~!/��|Tl�s
�g�lݗ���uL�I���`mU�2���)̐�2�W����f�@5�d���p7��=S��)����s��&�P>�atw{���mc�\L�gH/��f���ۢ�Aq��E�OʗD����ƿ?]d$|�������?R������Ow�Q����59�ɪN��]4
2�L�j�ɜ"�>��y����!�~������ƾOH�G�t�A�m��E�{�T��5�Pt����73�я}��2� >q!k̖�uoC�>s�2;��oVtE��	�mC�`��m `�G�pP<��h���	�<SpZ���.T����䵟x���D�}_��[�N�Rs����]Gu�v���xK�G�{Y8z>�x�@���>o�̡�um�uB��3|��B,��q,�Ept�lw
�&�e?����(J����\�M:�[�1�V_+������Z9y{8\���͒��:�JT��MH�\�=J���g)�d=Q	�sҪ�#�LC�D�@����(0��
ZճO�[�L�E� �}`ˍ��v�ǰ�jM$/R˟�K��������Q�w{�Fcٸ#b��fĹl۫JS8��.�#	V;�%����'\�fFQ���a2_4�.�s�3��sϷ`���s�����q����7#�K���<�S������)�,)7a���`ncNb��Ώ(Z����+�4$�T�X�Ⱦ�^�n$N�=��ד�D�6��(�(��ݖ� h�Ai^�dg�y��['�ՏJ�Ih�6��qu�ZoV"Bνd��ORBΥ�T�+���@����wn������{�?V�[?�h���� u9Z��ׂ����:B��uSJ�����}�:��6Td~�B|I��9"b�uO�?&�H��+�_��e
��*�ϯ9;�tT��ǀ�J��Q
��x{p��e�f�Vlj�8���>���=��(�#�j̉�Y��;mБa�$qa�+bRȚ+�Yԃ?���^����-��_�Z�ҕ�-���c-�q��+�����ZIco��<
x��
��1��2��K��!(���|utd>T�"����^v�)yЕ�h[n��(D�4��ʾ��T��Tn��s�M08	\/�ֹڃG+H ��:"���@j�s��<�n�C9��d��kR9�e�t
��w����f�	3�d`~#(�m����z�K�s�-�$=��{�OC�5�b�����ŝ;Bd$���H?lޘ�$��7L�+h�����z��������aNl�3_j�os����ٴ*�O��%?Vv'�0�<ڐ�l�C�(�ň��}������L� �g���Z	�o���l�?�R�c1:dհ���y$f������Q�xF .�ݐ�[��$�����uq�:�ǶR^�{<�d8���dFo�I�m�8z�4�R�:�׀���z������ۈ_+H�<>�k�$��EG`�YK��3��ӂ;�c��ܻ�j�Q�sd�6�⽷-˰=����Y|,i�?ۂu;'G7K��9n"rި[�nn
&^�� �EZ�����Lb� mt)(A��D��3���ʿrﰿ�a�ڴnM�kM�~i�k�Қ���IFH����TtarU34	%����(@�T�σ^��J���!�:bG���Ɏ�xhi�a��S�ԥ��0`\>�y��|Е�8��v��'����B�P�#Ϯ��L��0=F�|@Ydf�%X8(jIF	��+L�f$��$0urk�덠�sJ6{�S���E:�/��	��6W��yi@^~��<�u����V0fFyRE�X�PvY��[f���l��!2����b�>���pF=�g����V_�b��X;:H�z���u`q��z�J
��&v���C���!���a�k�l?������ہ�v�\��Cv �8��[9|z �n5��8�{iŅG�y���������`�VX�̌��	g&�2o�#BJ�Pܻ�k,F����������W�m�.��#R�Y�f�iK��Um���]����i���mY���S]�]|�?���֝&	:�vt��m`���U5Ǽ<.|�E$z�ji�Y�G>{k>�6��x[�5E��#�[^(�;d�Q�\��(���_m���	�t�����c/)�meSv�='����̤��1�E�L����|��	n�J�1��"&��֟Y(k=��h�a}-gT�O���\�-5�̹|]T �{��Y�LB0��5� �}}%�ߝ �6�>R�����CF���8�?~�̓4���/F~4�Ȍ'�bu�p��91�="H�q�ٕ�D��$�����6�s�1�l��ǥ���}w��� 2���D�	�hW`�8<�2��@ڰ�h f$Nm���%.�,"�W��+wé\{��$�s����>lX�o5RW��9�:�v�7��E��ϸ'c-\������������?@��p);�_��+�M�u9^�D#������~gʱ�^gt"7L%�R'���O���Y���H3�����*�
����.U.�s��������l���L�y;b
����0��N��+EC�n7�Wj��q�PO�g� EcԳD�<�MtZMID	l4x<I�n'��tÞY��R�CO$dks@�%��X&��1���e efN�Sh�_#c>�J�5���L��Z�~��e���(����22J���"�~A���4��d`�35��qX��~��˧ų���wF���=�?��k����FJ������$���73ˣ-�j�J��8��&�Zn�4w������o����(��`�?�֫jj��}�2J��$�t�j��7�7�Nȏ��Ż�+~/���m�|�0�d*B�:�g6�����E�}�,��Ό����{��ʊ�5�a9�T�I��OU3�rb3z׽ݗ�
ji|�ۧ\�6�\�O�R3t(�
uW��r�Z_[�}P�~Q�nb�h`�r�%}�����0	�����<�Y&I$
�����"c'JvRl���0��%�G�l�C9n��뻜8����R^����)���$r����-�>�d�u�,�5�wJ8����zv�P^���.�S��|w����敘0��D�[�^m�k�ݲ����~U:���=5�U����&9tb�8z�7Q�ĴN�������&�6���+{_{ؒ[��|d�ϕ��\�|$=���8�5-�ԑ}�tS�W�UH�z<��P�}�ߣ�-=6W?���G��ꡣX��I:S���|H�S�k�2����{z<�ⴝt�o@A ܽ�1��+�X������Q���!��A�)ô�z�Ph��q0�M��%�_cJF��}L�^Ϸp"��|�R`fjA���ǡA~OO�\��9��\@�U��tܶ�.�A p IpNsg� �[�3<��l� ��$Թ��iJp��l�u�~D�dmk�]
�ݭ9���^���B�w2������^�S
�S�C%j0Y�~�����y*mK���
K�7V���'����Jg��8�֙e�Mt�-)*�F�u31��*��󝹩��In�^��t�S{MJ{a�x��pϵ˨O��d���Af�|�Ij'�Yb��󧏼7�������x:��P���k��8w��
�%�
��DP=�G8���/��!mS���>���s��$}���8����a0�,���%P;+	�� �C;�a��E���Zj�},��p����aip��V��24����(��K��|�/������`������c����O��X6�ղ`��sC�ʩ��:]�����6*�\@�辠���#(��z�W��Śl��`��CBuse��vVyM'�fK׹��[�ҙ��t��Ȗ;}w��'�Ѿ��|�P�*o�r	#����u閈y^�+����Oaz��<|Z������y�$`�J1H3�^0>���\cf�ҵ�5��4�Y�b�*;:��|�[�t��IɎ�]]�������^�ʲqĦެ*G������Hy�(�s�t�],6̞�[��"��!B���j��d9l�����.���M������2�BP;�{���-�L��5�g�C�Ba�D]�_��S�n���[��#������R�W��©j���~C�3�w0��Z4V���Cr8A��g���r�|}��Q�������^���;��.I觯�8 ��|=�2G8ϸ��:��Au�g��o��5�_�y���h��ޢ�e�srr�b*���I�"�1&���ZH�,�Ża����h-�a�C�΃
n�c�|�->�zC.炝���QPH��5���̀-G��L��T ^@ٿ��d�D� ��t�B����-A�zV�����o�'����R�(0��B�k���ku�����嗛���׍���'��Ѹ�^J�'j��t�@�Ü�a��ΚY���us�z�!i�BFe9�nC�U�皊�9F�Dr��I�.���#�+.��B6��HceRd?i�<��"V.2B���%���IJ��z��c;H��A�C(���jxT���|*�����%�s��&�����+d��y���I�F��c1�$�>E��$ ��9��~j�G'��(1��,�G�6��j����~�S�5JDs�7W(�Ԓ,%�c��4}x�o��,W�-��9OpӤ:`���0�U�w����#·&fr5��M�����R������$�)�GC�@y��Bg��}�դQUW���r|�8�%��,t'�1>�h�H1n��^�e�ȫ�Χ���r_,����Ү�*������b*3	��z��$��q�H�y|��5v-�HB��e�4�ѦFC��W a�$ļI1����*��\D��[D�������l�;h����~K��6��}Dz�����u� 58�Fuܳi��U0����p�x�sX˶�6^rͱ�V���1<�]>JtF&  UM�k�[��n�"�l4y��ڬy���F}�/�zv���Cv����WBX�wc�6�&���ò����gD����\��Rpܚ��>���bf��/��YŇzT�m�D�-e]����l�<�,�'�t��� Aٓw��ne��Y��8��F%^ڸ�Lm1|�(O��ua�n������`��"�o@<㡈�3�����H��0t�\l�+2e�P	�UB�:�#7�yR�(*0u�M�H�@�T/�q*B�^���.ǲ%rMu_A�.�س��?f��	���>�A��(�Fhi���~.4BY1�O�'\�O��3U�5�Ia�{�ʮ�yX�u����-j+����?;��=祥���Q-�����%T��Ҍ<aղ7��+���]���������{��P�,K�������*�6V��=����z�j���͇�)X,O@�\M��aKE�+��ā��^;��GW��ΙE���s���)[��8����}�&:� Ou���p�|��N��nIb�r9:�;��`�����3����1���T�8��;���k�-`!��b��V
T�&�����V�֝����sS+did5;�ݞ�����P�S�a�H"�E6���Z�1H^���$��׍у�{���
x��[o�t���ۜ�.u����u�����B�˘1-)�	���p��g�hl�~!�~�S��
м�Ԑ��Y �)ZRȕ'p�Mr���XbN14���Y�v��V-Ě`&�N\��5BQ{'&��\�#�][�����h��ҙOB����c��,gغk�v��I�[��^Z�U�;c��h���툟Z�<�����.f���F�Mu!Y����q��v���Z+zkWG6�Ƈ���ǿ_��P��߬��!����f�ll�0,C��ؕ����_E�&:�-�bp�{�L�r_���b��.�ç�	�y�KS�ePɿ���@	�ڇ]LI�p(X���/ˬ���M�݅�K�|$�?1�M�/lHFn�&�

�0vQCtE�x�hs�֚���V|j,>�
�_�����K	d&{�GPTb.s���ወY4o�-�i�a�{����tr�f"/��2��RWK�/�l�++��]2���,�� E���obQ��]._�S �[�T1�@��O��dm����'��̙c��v���̡ NL���Ȥta�XeU��i��}�,C[ЫA#��7Yw��ԤDa,���e܎������KjY*�a{�z;���x2�uM�1!/�!k�3VK�ŏ���e����Iâ;�T	�/�t���^�`�YL�d��m÷��S2[�`����!�rDo&d���N�������~�X�}a������� ��I}S%A��n��_�Z:TE���S���҄���ס2�26�	'���V����8��쁛G�c����0����ֆ���٦��>��9�!CS�vy8�S�{@��&��i�B��ql��_9��3�}���;��j<�����������5�+�oRD�x�(0\@��g�:ؚ-��ey�q[
�\�3�����4u����7�[��e����}5�7����˂q�6�9ke)��e�t�n��Bu��2*7*⾗q@#�s̸��ވb��m�ڕ� ����{d\�UD��%HڳXQ����E\����]�;O�xw�!xo��Pm�K�!�x(�9솸�2L�l<�&0������D�6���B��Q�S��q��UZspmU�D�ʅd3#���h֒��0)W��� �o����[�#f�e%*R�}�|��_rl"�Zq�#;������ιk4Gا��,�92V,�_Y��8\�q�Kӛ�Ea���@�S�C�M�)������x�od��>�1<z��q������@����M,S._TTsGC���F����id�I�ߊ\?NP�b��@_��d'FcZv=%���Z��]��b_�Z2�6����,��N�D�\�
����]�����ox5V�� ���9a��������)������[a�����?�a�k�k�V�Kc�����M�}��Zܺ3Z�nK���z40�^�&�	=@����o&e.�����8iX)��%2i�O���=#�� I�)m�o�H+7�O�5�f��g��C�H�l��!�C�`�{�����+��3��.lh{�C��p��I�%��E�ټV �i&q%w��n�g_\�>��ƛ�\-���6F��ڶg�X�fpW^�>!x!�擘�.ƃ�����~�����?���0 �`Բ"�]����{eަ{:����@���݉,����o��$�ʊ|��&}��{|#���_�쩾�#v���=#�8���Rh!�r oN�V)S	��D�A�oIrK+ƴ@����~v\׀��k,o�Kw{��|�V&����Hx7L�s=Ծ�,&��Acs�3׳[��r�
/]s�����I��,�K.�cE��:1�<�Ru���t|�8�I�	S9ö,��+TFu���S�F�>:KĜ��M��( �|�$ܕ�'l^�Hs6�9;2I�πg�	+�>��|����	�\�},e/JZr~s3�;��}+LD�C����� B���a���+Xu,/�g�Y�_5к��|�Z=���ߘ�qtB�=��f3����Y@�����D�t�0P+�7�Z��Bp�y���I>`捎3�)9���mj���&b�o�qb8Z�Z����Ɨ�vr(���UA���H�Њųx8�/�t�4��{��z[���>פ&� 7
/�G"N$2#T�U�
�=N9�WIX<Lz�W�T�eYNN�X+d>VZ��}�/��m�Q���$�Ddv�j�_����\b�ɩ��Xh7�Y���S}+�1=+ ���-)4�6ț�Մ�k��U�� ��c;�Ԋ��þEy�@�h��N�Z��B��sP��EG�U������y�#�~[������/>DC��:�kP�m<�N�n��kt\\�+Q`��w��m�����6�;	F P�Z(
���F�i�đ�"mR!�k5���*
�
S 1�%�z�u�	Y�l�d�&��	�����3���D���i�����\�¤W���@��F���5��3;6?Ts��>���E|G��2�������~n�3���Κ�x��
ҕ�$�9T"FM�u�T{����PfRS;L��͓h����v�����W^l޻���X �����|URy�i� P�ݧ�aY��a��߆(�/�����E��j���ף����x�j����S������)o.�W���2ʹ�Ԏ�ʲد��"~��)Xy��6����y�c����Ԭ=�e�!�]B�_���S~��c�F�
'�uH��h��h�����)�j�����u!%�)zD��	H�_�5M�ز��ñxS�Gc >��];�%��澺���r�Lw���sc,��3��;�[�I{j�q$����oV�QO�8Q	g�������>����I>F���j�,îD�Y�,˞��{�<���qvC��O�z����|�;K�D�-�dc�=�q�z���1����mv�-�#X�B=x�Yg3�:�~���>����������0Խ��L��k��%3��o����"-5�I��4��U� p0���M3�D���V2�r�9����L�w�R�Y�ҏ!�~�Zgb���{��K~�$jA���3C��]l�X����7�%�n�P�ta�/!a�Q�q8��z)�q�H��2eÓ��.�l?=��5�A���O?[F1q��M׹K���|�6���qRj0H}0�!N@��aynP*���?6�Osp����s2S(��$��P�>���ӍI*s_���;���	e�Δ��6ӓ�&#^8�.�O��l� f�~��)Oc���H!����s�-:1�F�SI'	˝T"���?�n��;�f�%��݌۫g%'d	�L�M7%���!��0@NБu����Ί*���n3�j��2��<�5z�4���]q�x��hf2A=AY�?�A���:G7I����7]8�q��}R�(��7�+���@^���ʇ�{Dp�;��A��~�� t�=5Ш��fF����FZ1�xKB��ל�J8.5�)�u���
�+��Q���W%�����L �����'��+\Hz.����m2�Q5�@\��_�Dt�pA�3m��#&E��nf��p��M��lzB�L�eY+k��ϓ���)�����ne���o���W�� Ԉ�y�Dk�A��Π���V��u�ىI_ӷ��%����_JD�[�+�,�����շ�T�k��są�[p�;����])���4	�~��0wƆ�XX�ԺK��7|NxB�w-5�L�y�~���-�N�j�,B�a2<�ϹR^Y)�}\$~3��{/��X\9v����r�KS���5���p��X;�K�����4�Yץ��������1����il�!E7��Z`��9�S�3  ��D�$/�q�F<+�\Ap<$�gՅ��@Zf�~5O��)8�� @�b�=hZ{��<q�o�P��đ���"�hǋ�Poʯp�{��J�1�bF�WV/����<�����i��'1��11�P�{k���'�R�;=G��!S���\��D'h������{
�AY ���2�o�pp�Lz���2-�.5g���\đvfR��L�{����2��;a�;$f�[��ƫ̓RD��֨���t��pZ$�p��\��Ƨ����V6�k��]��1�yn��Z�l�3޶�Q�X`J�}����{x��{���Ӆ_����И��1u��j2Ӆ�=.őG ���b�׉��]��ظ�i&&R��՝̕�Z��V�բ�N�*l'�2�8���F��=���Y;4Os��R�[v8;�C6g�%�� X�@\1�v�pF����䐸�� =>����R����	��x�:\|@���7*�NG%�N����2{RQ	Bm-��$p�~��+��Ou	����%�`LY*
R���`Re��o5����x/��1m 4��?{����Y·8q,������U;�d�|N���Y�+��N�?b���/*�C���tx��ĺW��t�	��i�l��Arp��jm�6���1*�Sƞ��Fb4_宔4<��r ܟ��(A��_����U�����O��`�IM���^�HAݮ�����I�\��s�	�wZ�@݅�xg��!΁<���ݡ	�������t�nb�]Ql�r�����i+GK�:�6��Ê'ٌ��$9	h�Wi���z���9/���hRSծ��<��@�+����>�J_9W�J@V�nn���3���J�P{��?�M�����ט�m$`F��G���ۓ�	;��A�f�PW�{��GWC���\�x�rR��y��K���6`��	�I6g���Rҭi�Kd�+)�R��#������Eƻb������'�;�?�dF厜I���hP�[�H6���<y~u�m+�D��<�p�f��?Z��&j��НY�ӳ��o5e�[�8���s��i�ӻA}���[x#I��Zp�W��+̪ ���g����VG�����屺Vg����E��b�,�`/�Z�99ʪR+���oU�fSc��e,{Y�s�I���/��|�N�Z�ǻĺ9���[�L�_|rl#�|�_<��cH�s��9�3��ޫ�oR�!i ��tA���:���Bc��5n�	jI�$�y@2�軤Nj�Դ�D3�����$
�iV��F?J�)�[�٪��ՓX�7pO�f�B�h09k߲ЀkroNC���j�\�Y�S�U�(2��}P���鳘��쓓>��ܮ�L5��;=hu$�S��`_]:�M��f!$S���i2���b��"�O�����>e\B���(�z��i7�+0���f�z����s:ȃ���|���luq8@�� Q�b���q?��-޴R�VSTi��xM#���+�xl��7S�.ǜ^:fg��m�=i|�]D��O��iM_��@[ ��R� �cs?�f/��a�ˣ
ȸoq����d^�V�#�w�m���9w�ʡs:.�<�ͼE����V�L�m����uL�v�:q�(Zu�)}%;�Y�����H���A�e�w�?E�,H(�WX+����ȅ�O�86���6�k��[�Xw�Q/,�c~k�Нūh��C�ҿHR̄�d��������RWy�r�ώ���6�	�^�)$-����1TF7K���:s"S�u���l�6_#��#�XAJ��
(;�l[�D0E���l���N��``�z,@#Jݪֶ�'���*`tD$X���:t�H����V��n��&��8C[N�>�a�|�04P�J�NF����x�2 P��Fj�����]T.֐cw ��Noy��N�+��qϩd�59Yn
�/ױ0B�ށ`�_^`&� ��S�sdj��'s$n��d��O:�=Y��*��B��N�KQ-Ɋ�p�];=�ni=�qN�D-T�8w��h,����r� 1U,8� �>N�Ǭp�jF�1��&�A�X���=�VEz,�,����Ц��TdǸs���Jp�	Dzl��~��[�8�i�)��"�+�h[:���m͒��f�b����6��tm�x1�)]�,���e�L�G)M���@���X9���w(�$9��q^/a�["ݪ5QVO��wf�3�|���̃=��:�*�����V�p��-5Mƻ-M����5<;��*��s�#��E�˳V�5�Ӝ��|=���� 	��vc�^��[�
U�tHM�H��hmW{{��P� "���a�;��+���:J�x��}Ay�u'�>#3>�i=�2�&2�ߊ�ʬ_���3�'u���)���p�S���F?m	�ʌے\�5zov�O&.�~�X4��m�����2;�k>����U�p�RM�����z���I�xPQ@5�H�8�qt�7�(�F��к>	�z�eF��n���隷^���5o�$�2PW��ѥ'ԣ��g�#�{���&��֐��*�`��Ȟ�}�G�PG ���������� �_�+9�)X%�x�<ɘ���>9,�d��Q�0[f9��o��2��t"�]Z�Dd>{m����Ӓ���E�,:E�a�[�tDs�0�)��b-�.�F{	��ig
:���}����"�9���wK	��9\�j��([�لDF^�I��@w�Ô��E�R�,a�(@�s��G���]�|#�' [�Q)^����h�֪��E��p�=I~@DWӳ3?XP4k�o�̉*����W�ϰ��j�9��'�|N��H��,Ey�Ǫ��[�5�y�S��D�lv_�?�P�q[o�g!�=�m��ba/��y�E�rl�����6I�$�?���T�z��X�Z��{��%����"�F��L���C9X��C�M
bQ����8|�(�q���w���^mZ��h]��E4��̔��?J��>����f��e~b�m��}Y*U᰷��`�1�p����u��<���<F�P��"�����k��;�;�Y���֭��x���j��`<ta����>X7�N��@�Ǝ��Q���H����"��C�}b�4N��@ep>�<�%,*1�B�7R��\�q���-ڋu�O���y͚���&|M�9)�MO���죍�x����/|;/Z�eo�*i��0�}�A_ɚ�<������K\�3]��t���Cⷣ��{�Lژ��k�F����jro�#f�GC5�PDx����HYy��RrZ�0���Ef�.m`��!����1�{������v�	X��cq�w�Y_9�ܯ)?���3�p����E�{�Z$]�`Lq�'����������q2E��kDl�Y�_e��־n���4ba7�� ��$+k�	�]*�4FPy1C'y<�K˥	�y��rz��tu:{�������7�񯰻�� U��'�o�g��_ǒ90�#�7�k�m/r��$�J�����h
;jUdV�f1p,�=8��ӧh(��9!�,s��x0X>��M������/���>Ǡ=r��i��lo�w̧x,�!��خ���]�`�[S4W	���	��g�=�����F&�2�I&.��)� ��y[G�[�-�N2p�m{�B���c�!��`ȚbeN����+�O��K;&4�S(n-�9s�3ޟ[��5lK6����
��L=�czp��1�v�cE}�X�6��٢��lSW���l^�Q%�*"d
?�MO��</����	Uhg?_�_��	$��E���*,YK"F�H)��:Oz�L�`*��N��**5�@z���Rl0�2�c��w��/��A4�$<��SU	K!��a-��5Zk�w��q��D��j�A��d�v4r�"M������
�"�'���E��Ι��sAkcG�FG
L��O�~_4�d�ȕ�8�f�504�3�Ok�Tݾ�������"�mNj?:��d���N'Oh��4��7]�*�5L���[�Z�H:��P4����9��g?�?&�z�8`E��j�n�}�ar|}�|F0p+-��)0������3-�el_i	Ty;[C��R"U��ĉ_��ƹ�*G�[o�nvX���L�ʭ����d�^D`�tiW�!�N��p�Sx�<×�����@��
_z���ʽ�^�`qv���m��:��#���h�]̏hD�O?������k�[�0=�9��m�f0Nx��P"/�P��8/��n�5�1��U��;�pᵟ���I�s��	�����b)�D�@=[+�:zX�4����.�m���Z���b���S��]�ҸC����j䁣������xƵgi��������eR8t<���k�<�����;�#���Øw$�w���(F av��F%����ǝ��Ӫ�I8ֹ��r]�����j<萕9���'>�}���ź��\��=p�R�3����e(��b��5u�a���i?����n�-�S�"3�"6PH���|x��q��X���5<��*zB��Mw:�R���1s���RU�JW}��������{�.�Vle���{"��V�TR�=$�o��`<�J�/oN�]�0�(����w��������G%���d�C�*[�̢k���^gu~�j�������so�MH�읪^ᅢ�M� ��#�4������38��;��1��-�t)��:]4��߬-� ������-{�ޕ�a^�?]'@��yQ����{�Hy�/a��}	F0�8!��{\q� ��!�3�a��� �%t�OisM�Ѫ�;��fh&����wc�\�V�R��}��k!�N�����a��ͨ��Л�`O*R�Ia�8[/��P`��,=�}ܰ���o��`*̳�a�"iYw\�^F;���4��.k�]�YNB���:�!{��~�ӾLk�E���V���1೿)�xɠFUAPg *�Ѝ��z�l<'_��*��{=�K�ֻ<�B�r凚/�H�09��=U?��w�s����w3�����4��>�ǘR�����w���ܜQ����3�M�S���忻�C��3���1/�����Z�1a�y~N�P�pn�t�<�F5sp/΍���2��m}J�Jp�A���s!@�8���k3a�g��{��/7Y�ϧ_�5$��G��N�N\;8ƒ���'�n6��`E8�ĭ���k��{5��E�mY��H
����~� �5f���DXD$�=P8���_�d���׻
s��KL+�rXo�n@�~h��5/�w_�kP��U!�6��מ���ߢ].��G�q"(8��^�gvS��Ǒ��SC4!+�C���p1��H���'xj�ެ��9�Oq��f0���������|G{�v���Sy<�_~m�6��vv���L���":����_w��O�s���"���@,�yo�T(��_�
*�fp*�:��+�4��IV~�z]�rՈ�,�S�NRZ��Q��͖*�Z����%rN��S���NLz�B����5'�,m�+�"��Y���\C��;�Ik���^�r��|�^���
��ɉy�� �y��y��yПc���n
Wa��,y�ɿJnW�an�G7��ܲB��^d��0�Eۻy�)�:��i0�qǧV���ʪ����b����Fp���cu�~ߣ+��T�G����f����ҷ�v��
S΋?]�پYj��d)��N�i��[ԱҾT]<�p]���9գٕZ��{�L}HPg]D=HΏы�����m� �UǔTG(f,���@��4��.�����)ў�z�׊pC򧥿�F�@��h�4��/� ͸5�\�r%��~VHR���y��I8�Zk��f���7Ɏ��iF��S���ZT�")�%�����F�T�sdD\���[���ť�mIÀZ�L�t�Ǻ���;k+`R������0)��Ĵ(� ����~]�_Udt�b�KHF� �>Y���e3��M�^ �R^�U|/>j��%�tFR�t�kw�#�s?u"�94�PSGm%��p2ٹ�W����m��R�a��������v�'���@�6m��rj4m�pz���f��J��E��6�PZ+c�յ�R\�a�P�LI�����_��n� �
ߦ��w�m�*s;��� ���7��yZ�ɐn���Rl ���ID�S��#J���$��
��gcԼG�L{��E89h$�F$a$t�tX��!�]�:��1�L̲`m���Bߨ����B��2"�?[}�CF�,�}jYBλ�I�&�\�O��D��)��X������t�6�ΠĨ�Q����V+��e;09���!�y�dK����g${�&h/�Ro0�f���P�^�����t姶���N��Myw������P��o�'ss�G��G�I��`�TQ��������l2��-i�;�)6���VH��Avp���8�yi*�͡j���EIG�<N���3O�Sv�l׽i��!�Q���H���65�Aj�	������� �.p���*�ӎQe�V�)�jXc����q�ɛ���9�'O�8�f�_@w��NN��Ӭ����%�}�G�{HX�(��Tl�D^���P6��7E�"��~%-�=�]��&]lsq�����g�i(�P�t��eK��?F�L��f����!�4s���Ҝӻ�29���7���gF��L���d]��FS8���ci��9�<��0��#��(�~�G��k�`�G��O��%��K�yE¥aI$b	�ݧ�yd|�Y�'zQ��E���Rt�]�HǤ�3�֓��ߖx����p�k�!�o�b�����Ho�M��xԡ!209܉���`i��b���dɝC����^�`�_�v��a����9`8�:��Y�;<z3�bQiUK�C�����;����""jU���]��,S��Ap���(/j����$}�s�4���l�K�d�ڣ�Kk�+�D�}4ņ������T��^�#�)����/�$��_�:�/�Q��#��}�&�0W���;�&cg�<�w{���*(����.���֝4qfs(R���Oo 1T�J�c���+T�ӜV�&�u]kP���T�q�P�,�S�A�j��:н��[�u��_e�Ac)�L�іj2?Ԟ��*d��n�S�:lw+3A�,@��AGJ���H^�?F���Y��.��Ea�X��1=�c"�!+�2�e��dV��~�]�p�(�Y�:�{��1��>2�9-��ȗrKU;��A�A���(���2�"K�������+�f�$�ʑ(������J4Z*~�����:g��m}�M8Q.{��4�8�$�����2�>�ݍȎ��W�u rLp�JJ�|3�4[~6dtx̳��.|��[�YB�׈٥��$[JNuWJ��f�
,x=���)}�{�YoJ��R�N}��Xu�ϛC,�K`��A�g�ٝ��t<P%��_��|�C��둇#!K�uY蕿,p:pB�:�E5��_�e+��B>,`��k\�J�[@+�}:!3-�<�S��~��'�Ż.T.Z,�D�=�%��RƑ��G�duO�N�ҡ�T��tpFT�]�ݒ��/��36���S������4�麼k�i�3��Lj��ԨI�gTG�(�*�F����+�&��4u�	�s
Zp\c���V0"�#�X�3�<��ڗ��@��>��B�^� F�H����uL�bpe]X$P|���y�v3����d1���d��v�	��'8��0>Ā��J�I^�JFߊ��B�m���.��1�bt���i��'=�� Q�H�nlW'��X�I�З�ނF2��j^��.0�u1����\�@�YD�2&�z!SHh���%	ʋ�/�_ͪ�h�)�N������fD�4��mj<��=�cV>�	k�{L�K�߸� 7� �oH�/ĉΌ�����➡��A<'�E�=1Z]uH*9ݤ�"�~�gL@�q���ֈ2|���O����	st�[z⧠N�WN^����42�5^�X���0xw���q��v?$ռ��Mh�/�o��xx�`�����p���+*��s���>���|����}��Yr�m.̀zDZԂ]׾����
;~�#ܾ/�p1,�:[x7��	��>�_ˠ�P|w�G�լ凌�0���ߏP�j�A�_�2ew�Tebr[���L6Hc�mî���f���2�2`��o��Ӯ��q��L.���HT,���X-����}���������ч���hYk�N�Y��n��K�ن��n�$�22��q�
c� ��PQ���R���	p�����a���( ��
����l�||]f��N��q͌����	-ca��+����+���7�edn.�*g-u�[ 6)t�_#Q>y.��0 ��q-P_�zߙE��b@��2�}�s��UHR0��Y�H�� ?������N[ua�<�:YF�Uxӛ7׃�M5Ԇm��?�B�)�tu��ׂ_��܊�o*����l���>��� G���90�*u�&�J��DQ]�X~Y��_\u�9l��Ak6�e�9��D����+�������z�qYH�,�z*�)zH&�1�8ٗg����c8�.X���Bt{V�.������C���*�Q1FW�8p���6W�����ǀO�m��b��x�����������t~l�!�Q9Yw˥����5+�b%�Z���t��܃�Wz>�#�(z�����k$i�۹����]��(�6'$��Ux���b���Z�����#q�b����($��W���J4��m�1�aT�l�Zb���fR��	��3CSI�y��2.Z���}��{+�a�&���D�~W�>�J��W�쫿�D �B���G��ky�\6z�mB��JI?��;:��2k�Vʊ�o�r�Aa�b�d���fNxa�¿�Nd�3+m/�Z�!�JU��|�6�$�w%��Xtc�����S����TI����--*�?)S�6�����z,�3
�X'�:�,�>��V�-V+Ⱦ�"]ڱ�Zߘ8�������eW��ï��8���-� V7\��4y��ۘ�k���Xb����)�D�6���^��eZ$Mi�#��oܙ3��w9�+�Ya-/��k n��]��jh��(��v���F��>hy���+_I�c���!�5�����wU
]t�n?�xT�  �h.G7�i����Ɗ���@A�?�&����ր؊B���WX��	j�V9�DaeA	�9zv�'���f�����l�}+�Ľ�~b�n������3��K�j��E������:�P�|aDna�P���=U�O���11��<��2���YԒ(C�����{��h/�Q��#���;�/O"�K0�3O�p 	���x1 ��9��:N���]z_�VJJ���c���[�!�X1�A�TmJk��I���@�����>�E<�n�G׊� G��(�?t����I��4A?����?^�P��� ��<_�c]sUb�����O���c6g�DA�U۱�]�[���2�������<��>�����K�Mȃ��95U6ɓ'�����:�Ee���,�jd�R:��b�`U�ǎ���uJQb!��qK��� ѽ*9�X� eB(~5��~/�y�Z�kU8;�Q
~I����-��x<��!{�u}i����N��І�ɡbNn^��+ΧHˈS�|�ᕃ�-�H�h�7�ʣ,9���hE��R?N���,��!?�W�U*��zI/��HT����$.��	�*O<�C�֡��U�3泎ɴ	�y!j�
1�\G�+{�?��.��@���j0_j��3�̛�a�Z"hõU,̤1�)ƈ��7�����U�	���\���e�ϯa�ᣵ�/�Up�=�kC���7ߟ�7��) =��O�l�h���
Tsb�)}�R��Z�澣;��ȱ��= �s����9��m����x)	���y��8�3���EA��y����E���|���{���7���_�ZW��3�ӟ3�C��P�M���_�����������d��Fd��V˙�|Y�Z-<�$��c��t�$�.>����D�\��/F��_#KK$��@�+fj�a�AQ�6���>TAdo�	����4c ��/?�z�DH�N�:R ҦgQM�QK�����E}�nf��>��M�F0�]D���\�n{�sZ���ʳЩ�<�Nz絾�x� �vHv0���y����KKL�0��(��C
4$Q����(\�uډ�h?K�
�-��І�e�m�����i���7a��t�|P�\�gI	*��V�o�	eX�ՐFA�R��x��$ן��C��(\,^���hg��+֛���/�P�+�bޫ�d��F����K˨�4`��y��k����&Z��1͢.�ws2H��Ǧh��sBJ����6ܕI���}.�1ı[,ώ5U�X(�� ���D�Ĭ	i�h�; 뗴�я�틗��i��l�	Q0f�����<�T=>)E?�\4����u�/	<v�=e���*- �C�>�ڨ�`�M�p5���g�C������@(�IG���N�oC�țn<��LY��\��T� ��S�,jv9�����Lo��6�!�tGx	$s6�q��@`�Vpe�T_�Y��{����TS�S��UHT��	�&���n��>���4\��R��z��-��uփl�x��3�Z��To�3��7}�ׄ�&���L��o�1�v�~1^x�_�Ax'�sï���j���ůOV0Z��|������.[�׊t���������&�"���!�yy	��1}�n�S��n�  �k�]�����fC ?�$��ߏ�l�ߥ0O-��rۏg^0+3�����m:L��(医b��E�}@��]�_�M�c38I0}cB@6�A���N�\���!���upX�o�J��di�P��]�����ѕω�l�O��(��y^�*����Գb�$RB�ТM��w��;�>GN�4�������q]c��&0ԃ�c��o����m_~R��t5rʩd�tKz��Fn)�Z^�$m�'��+=�*#��SJ:�dP�C���x�JܲQGU�ҬJ
�9`�a�R�ϯ+;��(�e�� �X+�}��z� ;�c�p�(c�F��'̀�?����k��i#�a�e�\B��l�����sS[5_��!�z�0�x3��kdKe���;�ZTudI��<��,d��JO�������@��� �	2�klX=+��ҘOT��/-�������(X�^�N\Br�2fhx������~�-�F,<�F�62�6m��X�Y6p��(�<��NG��g�3k��P刼��.�]�8
�����0d�t$N��i,I*RQQh>��*�R�4��箉�G'�<�� z�2QK{N�o�-u�C@�ɭ�a����� l��J6H���Q6�(@J~>��|�F(W�*C�BT��������AHG�2�j�tV^��i:4��t:����ޯ��`�`XR�:3D���UBn��Y�J���"�O�/��|B�'��/����=1>Ǖ�\h�ܗ��4���Ţ�P���W�N�D�~ܫ��&[;��S�gXl#Du#�ڭ%z�V�u��f��y�,7!�I�]i֨���1k"���0��寁%Z;7��u("'B�u�X?w'ɶ�,����c�B�ALN�n��]���1F!�	b9����`P�_��4���!  �А狫���׶�łNP�e7�[:b���V����G~}�L����>�|�jZ��H�ͮ��N̅��r��/�l�qw�J��$��׺�G�>�$� F�x�y�aL�h^w�MC0� ��m�h��j���+���p�[��K_�9 _����� W�\$U�`>���To�j���zA��F�6��V
l��?�m�r�@���jg8x��H�bަ�@�W2��۳)A����Ώ2����G	xo��;�����xi���~e�����֒��H@����.h��6v��W�.��\q-�4�GAM�wS��֓PnιV�(���]0���� }�V����K��o�EP�~��T���IAɜ������Pֻ'��maԐ���|����n��a�l�o��]�8��.�|��Z�� W���^"_�_��s?���	np7��#P�>1�Ku�k�T�"�5P{���3�,ˀ<I�W��O,W��8��i[Wt���vjŗb�o����u��A�:�9b�t�v
��.r_h���8����_4��E��ިGٌ�ٛ��m*.�]O�G�Y���
F����[�2���L��ę�b�W�5M��)�I ��|�oꂪGt�7i{U��@24eZ:�����/�59�P����N�}�x� ����t�2h�0���D~�sAJ�⮳>/(��m�u���:���{[V������G>���Y4wUML�yfR�	�I{�����<�2����T�90^�������
���F����<Ǳ��"��<�[~k�a]I�S]�A�}��<�q�O�?�ˇxB����嶘����jy�Z{��es庆���T�C�Ha� ���g���Z�">��Z���mG���۰J}�L�AVeDt�&%�QC�W�&��r_x�	��L:E��(\��v�}qN��'��؎�;��m�^��6BK�� 3��(16]�^��
���:a��gQA�/=7��[L��k�-Tk
|5������{qs�ݵ�.��Ey��]kÚ0�Ԝ�c�68��_�-�ˍ`���^tP�)�V��vD�$�5n�<<��q>�����iL,*���71pu7���8�V��g�,�-1_j*12W�G.��»����)��+�ܫy�zz�sRx=����*u2  }�ɺdYo��{#t��CZ{
g�j��M����G!mJq�Ź���L����f�#&����@vN)F�m_�}n��)f_��=>G2w�P)A�i��G��GŀD[����=̲�����f,=A����}SV7O�嵆�"e|�[����^��@�~��-�.���y��΃F��ؚZ���Y%]nSd��-6�;��;��>��%2y����m~�zc�fHkϤ\[���x�K8'�tHh�[[�;���>%��5=>�<�����\��o����	:-����d<fl��r�NBe� iW����|����3��}	��E�N��a>�]����g*&���e�?jlW��
��*P�^@~�q.[��>��� �kNe�ӄ�����I)�|O:����G�v�P�G:`�j�]���N�$�� n��i�����TEî���<��|%�@)�M������r��B�u�R��,���Uv��aJ��t�	śr��>\�t�@�.`l�&
�(`�껻�kDj��oȗ���k%rVkw�4���v!�G��I�7����O � R��t代�Մa��qԚi�%qZcGO�ĩ4O������?d���=3Z�f����EN@��pL�f��yڤw�Z�Ä\;�]�.f�B����U�D���)��W_��lQV�#��LO`���z �P�E�������2u�F�{�rJ�F-�"~�s�,2���~u4�/�;�'�%�M�!�dx��t�4B����=?�c�z��C�������m��X1W��D��)j�1z�?��B�[�*�����םd��L�U��`�(������1� �W���ٸ�B��+�(O���=+pΈ�#��Y��-"ZrF	�e��y����d;L�$PtZ^�؋5t��8P��%.̀1heU�i�2״��Ո�s�'�qqO���B�j�㥠颿�~Hg����F�b%{��Xw��Wn`�7�֨y�c�u�o�8d����F�����۹�d ������d��2b,�^L�:Uz��6��u2�64�$���F�ir�Y_�퉄+ѭ�n�t�l����g���0�=�R��ۄC���0\�Dt��ɭ�V|ؕj2zl�|qU�$���M��-�Ihz}�a� d��e����g��|nA��{F��|����
Gã�,*_�����1qTQ@���hX��Wt��[�y�n/nU��e 4�zS����*r��=��R_2�w��[9';�L,���Ŋ.X�͞�=	�\\rf��M�L�L�K��SX�u���=3R7��1���j�Q��^���ݑ��/�Y-��!Ņ ��o:*��Է]�%㦾��W%����{����Yi�]q<��8N� ���D#��KѴf}I{��8����aݞg����~෡��)�J"�+�\��4��1���y�+���~�������+ޛ���#�����sJv��4�����2u�9x��Zh��*Y����]�z�3YO��t�Q��nkFѦ�g�gb7_��x�v<%r)�T�H8�Q~aw�l8�ߍ�9I��E��f�s�#�Nnv����b
M+!���Q�)僜�:ǐ ub�]x4�d�Oa���52` !��g�"�p��{m�rTj1���Kl�{��_C�5�$�ÕH�<m�J�_)|7i	D��җP�|!$n����՘��F�O��˦�m?��0���?� 0y\���L�;����r�T:�/>�t�zm�B��f�ۤ�x��q8|��Y<��������ˊk�U\$���*F�Q����	�5�6r�6��Ӟ������ׇ�
1ՠg�JC�c?�����b�#�Za�����_�ΫjCֵ46�a]�%C�n�>I�9�C����b=��ϗC6�iڼ��X7epZ����3���w�4�b���>������u��������Ң��)���^�C�-V�S�
��/���Ţ;����n�"�%�o�,���Ln���  s�[��H5����UI�����s�DDM��N����7�cP�ѾU�#�V^6	@Pt��Ƃ^w����L��.ܶ3�A3�f�����ƭzS:th��1�j����6i.�Ö��ɔ�Sw�^^Ȍ�H<%T�~��2V��<��jȻoN�KJ��_��;�����^K-�1�K��N+����P���)Ks5W�u!mkU�1Q��a|�dat �<���V�w�
ӈ��nT������/���ʜw��l�n��H�k�<X���s���?�X��ˬ���������r�jk�Q�Sr7\@+0�)��mW?�[�O��@�q!�R(��5?ݶ+���r ϼUw�6�f7���ÏŅ� �<�S�>Oi}�7	`>�3A�P4��I�]
�d���+����(�h�s:����#M��>�̺�I@-��1<�:����4���@��;��$�����B��iJ��:u���=]�`\��O;=�{�k���ԚaI��2|��n㪌�~̂�����4�4O�l ��	�ۭ��+ݓf���dK��P��
c8�)'0�Y8E�l���c�J��������V�Cr$�G�c�+�'���z�7�-ʝc؄�Ͽ,����˧�J�}a��kJ��$Gpa��P�����q��ŧ�:�����*`H��{�wv��-.ƅ>�2PY��/��W5��7+�CF�$�E
ԉ.
�#������	i�� ]��,�}�jL�BeV�+Nj������e�b��]I����3aQ�A�y�>S2^�+�l�m�$��y\@fA:ŵ�H�,�gQPdX��E���xK����	�/�5�9>���m�!1g��6_�zˌd�M_�A2�`HS}¨H�����]	�3mS��!�Ys3��I��k���:p).�l���GY���{f"�!2X�k��H�� �'I�{x�,L�V��ZQO�O|F������؅|i�^��?��N���Ή��K�CB���S)z��v�o�xS�
��))��o�G�� <��b�Ę���9��)|/�N-_t�(��i��F���)o��nb�,v��<g�9��������gD@|S�1�[��R.���Đ�^�AYנ�c%z��ݠ��|vM�t�J�౛��9C��;'�v F���5��+߳�}��h�&�
8�u�كSn���(�B�5~{U3"he&F�*skͣ��K)��q:�iE�SS �:�'Z�γ�A�蔉
=?ZJ,K�ި�(Η�P�OiLԞ�M�҇�AlzQ	~�gŪT���V� �j�J�y(�˲�|�o�g=��ƵC?Ly���s0���%ZWr�(W�_�%Kx���r���ɡo�|f�8��yy<�Htx��.�]�ꮦF��z���*ba�)��Y�q�)�3�VfZ���'�8��e�o�r�+byV3~ABձvC5�(�yٶ~ F���y��Q1�J�h�
`G��_��28s_����������16���4BЯp�h�"pz�8�V"'S���)6.�&uQ����r���r��'�:��ט?�U�g�j��ӔF���M[E�=c�
!:��٣'��������F�XD���(�bL������9��@:���~������;��Z�RLeKw���C"��#Z���B�KJ�'�#�?f�%�Oɇܺ�{��9>l�1��vx%xq����K��+*h�b����gs����]Oh:�F�.��!d��~tڳ�a� J���V|S�?\�/;H�4���,͠�B�8lr/m�������u��~�A�0!�HV��	ÙHݰ�?��X��x��"��aԌ���(�a.��H���o#2���+C��v��KZ�"�RP��T7�i��-���bg�AR�^���e�Fl�e#eKT��[sv���țni־ |�b�<`�y����%�S2���~g[�QOi�?��>y3@��*���y�Ze��&څ,�鱑v����w�<�e<�	�X���h4�sůQ���Bxa�1�U�L�"�<~�G�t"��Cr)��p�-\��֤��/tie�`aKg2k��?1�"�o� �[Ts�	7�80��n�\�P�t��Os�t�w��L&ف@ڋ�w�Y�c��F��s�A���kC�8�6���+��^k+S���x�a���t�'��V���y���<N�_%H������+qf�&��Y�wcZ�a���:wgX��������������5;��<ad�"��l������I���~%$p�u���E�p��w��I�k���Dxj�Q8���l#+1�\�C�rC��T,��bL�&+Pgpq�����8l���E�]�^��|����.Wu���I�e9|e>@�`�
�\.q ��<6�dW�C�H��Jf�k��o7�j�%�[�z��Z
d����a(�?h�4X7�Q�*��n;oc:&��/�8Ck�Յ�bb��/�������[���d� �y�������9����+]���5��LEE�w<W��{JgI�������鑆����ǀ�����Rk�i�ٓm zNG,`��V�u���S�3�)����|>�
��5��s*�"͝X��5�7}�0�@�F>6t9�`IIYXI�F�J)8�"oO����($�X������6F���������p~j���fk���/�@m�G��g>8���H�a���sl�4�Z	�����J�5�~��H�E�����V��u\R�L�[ұ�� ��0���"5���`-�O��޾tPE�띯���*do�)�q�]	W��x78����Ãu����Ct�iT�4ai�3p6��A'�8��G�"�V�d{?��X2^����Ҟ�^G�\�j��Z��|*� �r�`�(Vj�Y(sA�ϙ�	��jU]{MWK��)d:��p�V��cGU�#|I��j~a����}����W�!����s�I����4~�uUl. ��@7[�=f!�[xx���j����&I@�:�I �M��dS���q0:�*X�����'�B�O��s2u2)�o]k_
T7>hq�:erٜ�sp�t:2����#h$�Tn��,�^|MK�拫�n�?�rݽo���68�1�����IL���t� г�w�Z(������ʍ�j���3��C���?�q8�9�cvys�������_��XWRڌ���'���χ9\��'f����T��ݜ�|��#.���
��u�+4���N0#�Yip��~U0ٔ2�4�0=q��V��h��.�!�E��Z�vv�W�		�V��-��z+X�*���+��Om���w��6�[�e��4̩�۳.�����g���L�֎�a�4�b��E"n�U
6EuQA�iQ7�ɍ�)���� Ɛ���.��!7	2&�H�e�@�#W �辻sqD�E����;��|V��x1
�6u5���. ٴ�c��=�$׺������+��pғ����n�JϙL��v�~9�.���pHѬ���N���5��d�	���Qtf+��)yG4.G�2��E$��e�z x�ٲ�[jRϽ)f2��j�1s	�q�J{��Zi2�D,9��}���ט.p�X�:�Z(�VYCG�
������,;Y��үTY�K�O7�\��m4�,��[�0�l�y�Go�:T�P�
73��V +��+��
�8�cb��P�e���1�m�_���s�� @�Ie�?4��N����$_Eɒr�K�:�9�W26�
=�! ��n�����C�J��ɱ�Çǈ֧���rH��K���P�1�Q?%�
��Kg}c7;��BI�����apg���a+�əԪ�� ��.�l1�yo��pS�XzCa�W0^g�iN`�`�I��I�?NS����7������p�\�u���L*߸9)ɞx2����G����g"��u[>�^�bM�EN$)ً!���F��
и��(�p�#������mI�{�Z1v�0��r!Ӑ���`C���L�Qu�d�B�����A�5-΍L����2����ԟ��ƴzb�9c�7�,�D�qb����g��9/h�K�g-K����~�&*�W�s@@d-�nxU�Z�6/D��!���b�y�p:�S>����q��@]ұ�\�:�}�B��U���#6��}�:�uZ�ꏯ������9I��{2�����j[G���ن�����/���$q�4]�Ä���ÿ.�?d��D��(�vő�Rg�^�S;�<N�Tm�j�ꠀ�<�\2%]�e[jK�����$G���#��7��4�k�:K$��D�Ҙ�Ɛ����gpJ���t8g�LctsL,q3��?��eU*����l:i���+-Ǔ)�Ym8���/�A5|ow���� Cv�?�|.�(�1b�-������g��I8�p��:�]���XT"&�]�v�x� �M�����i�mj{tn���<���l�]uZ;Z��2(�>_oO��M��@�q�����њ' 3�/�=/O�h��Z�2D+}�f���g�Y�J�k�P��m+*�<*c�Rb���3��g0����x�;7��<�\.�lܤ �:�![����}����urL4g!�'�P���N4�i�b����C�mkv���@��h���@�@1�`U������J
�3�HlDb���WG��"�B~ߨ��b���m��Y�
��ُ��ؕ�sq��-q��LW��R �=ou�'\���O�r������N��#�E�K���k����VL�����ԏBc���E���%����ړ)�8�T��%������@�4T�����3-�1Ũ��ckL(O����BkYՓ����}�zO�A���/����f}uE�g�W�
4�2&��\��zt��N�RƚZ\h��:��s�� �1	?�g|��jM�%�P�g8!2O��͜��6Hks�y3z#��x`���%�Dp��Q�'д C��#���e��ԖaOe����Y�J|&�8p�$m���\�@��q׼�}��b�BW��.�0��\+P� 0_�ǳY��gO��ЋR��+St�>j�G@���
��پ Vq�����V���@�1��>�w��e�͂�-�h�ϻP,N`8�9������$�k�pq}/y	<�T!*����P�ٝ�Ii���4�_ Ƴw��H�'��X#�`��ēW+�M�-�rV?W����9A�� X�a��T�p�)?�n�	���S�V�`/�8�ў�B(�T#	��Gb	���K@ȗ�(�
�8�Ԓ:q�pu�aDI8�?@*����ӫDy8�Üً����	�&���{ܔ�M퇤�n��|I��h�)Q���k���5VjZ8z
�ǰ����OL��<�)�g3cԣ[���f���-5
h0`���q�~��Wr�-���xG�S��̲GL�-�88��drn ���/�:=n�(.=�`4�$Jl\�,�_���%c����~m���� ��&���ud�D�ta#r(�Ǘ'�-������=*�D���,M�s$����;���شˎ�]����I*ݽ�=�''[�}�>|a;�Lbx��I����z����'��Va��`�Fw	q�¹��&��J�<�dSGw�u� M-���x�wxQe��HU2�|��7�Z>_}��"(f�����N|�V��9f3��L���&�Uw����鞌���S�]����o�J�+]]ϩ�a�(¤sd�{x��%atn�*Ze���#}y��/)�-��X+�
��VzJ���X}v]Y���HZH?���U���}|��a����J�Єu2�ړe�eA/!^�˕m �����^sI��6��-�4]�抹&��д	a��I�Û��8�YQ#��_o-{�װA��z��=��jN#V�ݡqr$���&~C`��=�3��|��w�W{fx�*���{�3���O�	�0HFGl��^[﩯�jR{3�=��1Q�M���*AH9����c��:�;�(���������W��.�8�d��⑹����
*^��P]\�YRW[ ���P! ��\���T{JS�ǅ%�)"	C��E�E��R&��B���~^��t���lղ�G�xH��Ƹ�a)���h[�������v������kq�B�G)�#����8ޑĮ�<(k?~��Mn�R�8Y'��Ԩ��^[�|t�ޝH �~���u���6�?ٓ,�q1>�|^VK}=�P��y�w�N~'?b�/K���)�m1������-ߴ$v�B�#�E�0:�v�5Ȫx>���a��!������]�uM{��˔a�̙��$'���#��g�@s^�i�
�*�k�/�:�U=21�l��wt8�c���ZR���IQm!-YVN&2_�bt��)9M&����n�%���;2"$/������y�V��A
�z{k��'�� _:��U����e�'�RF�$�7�U�#�̐����^���ub��Rӿ�W{��Z�|�7fv���ѩ79�p�}^Nr?�mϾH��)�fH���J�f+\�͖e�Y�C�ȓ�.
�d|( ��!>�����n�G
zˇ�3�K�_����k�c����~1�Z�_ΉQ���\����v�dXi��F���<1��p���Ԃ��o��9b`����"JrI`�A��^�»����0)����6`g*9�?�+\B]RmoN}��+���@z���k�
����I�(��q1p�%������٣�"ײ��Oĺ�j�kCu��u1�����*6��V���-ޠ]69b��k��ԜCje��4O�W���A��f�R^}��MJA5��=;�ϴ��8����@�h��"���/W���Ml��M�#>I��?�e3� V�i���޾����B�A�--l ��$��)GkvG��/[���g.љ��C�v7g�e�z�(v�K�����Pa�Q��5Pt�ö0�i`L=M�i�� Ә�?���uHJi�`����I�3�Ih�t�]�{!������%W�D�E8t!��ƇW�!����@�p.�e ��w�X�"4%'=@�%hTa�ձ���L��\GU �ϧ��w�������B¬(��ѵ���·2 A���o���QTk1/����l1'���2�ғP`�?��*��&OŲ�K�2�T|B�OF����O��v���戼t�q�>h�*�@��<�+���y�dz������>�?�z�Ʉ��\-��ғ�Ul�'
�J���E�(��u���������=�b��(�XQ�}��F�/P�{`)	%u0��e���1`���P�sJf��7�2/�+d�6}��g���|J�Q6NÉ�%M=���ENj?���]�S��zDW�4i�@I(�s@d=��	 ��+�G���؏WEf4��D�L�� �&qs[n�	t�/�Uf� �USE8�u^�*P�+@��Ƿ.�S$t�b�?�Ȑ��5���ٽg��IN���1nt,��̲r�<�k����!Jw��c���@e�����5��X�y��|�Q�e�ږ )hB���Jѱ @kv�[<�b�d�
n�iU6v	H�M�{����)L����N`�81Y��y���x?:��?{8���ޛ*�F~ܣgb�S�qq*���*��nWv�ryy�N�
���jQխлf/'��~�5^��UFu�+�O5'��(�EI5�i���x�,�0����Тd࣠ŋ���	�>��("��Rx�fs�;PG��`��J0���N��sg��m�����3�1�:e(��d���x�,x����f��S��s�RN��]�l�<��9ইCɿMTXJ�>[v��,�騿���;@·���~-�
��Ck�ݍD��,x��|�ǰBW:����$J4������M	������c�,2�ƾ[�+��.���ڔK�|m�Q\N$6h�($r�/��`;�p��D=wPڃ�I��W��<��o�ۻ�x�u�%�w2�r���n�dm�Q-:� :�B^��������o�����aL�}����Ł�:ǈh�M��˹ƓemzC�p|�eW�t�v��x��Zm�<�;o)	o\���VG�����$AC�x�5��F��y��#:��>%r#�e$������,��6��y��D�xy*eһ1wէy�
���� �������4BP�qA�
�e�����x�[Z���`�v��]�W�C�[y��6�0��d�V����fHr`��p�#����LI��
���N���~�_\?e9֋I��KVݍ��pb$�f�����CรP�暀�kSg�G����gl�ͫ�ҡI��jc(aL�V�`���i��b�ʌybV��Z#	��h���?Z�x͢�ۓ�J���Om��4Eq��)0h��'�T��er��&2f�G�ݞ��U���ڒ���)ޕ��'�V,c�,�x�+�	�[T[U���Y��G��"7l�c�;#���i��s˪,J3�r@����j�MA�"��3��"OW�d�i� ]�K2@I8�fXv���K���[e�mCq
]r�y��40�O�!��Dw��ǅ�����m���Ē4�72�2�b�A��J�tz�����ĉ5����3e��W������i���_�ko΃����Ã���U���T�tI�4uP�O����{���!!�+̪�d� *1�?M�c���~��9Ӹ~�(l�A�~��e���J��I����}�����4e��:��X=�3��R�f��ӕ��2	; M��MdcDY���Z�fчJ~����21o�f����ŷ��8��X��|m�����|J�z���_�䬔t�`.�a2%��@H2�5�JC�[�k�`4��U���%݄�r�d#����;�'�M��-�潅��C�4�6t���=�����?��t�&�mF��������b�7����8AT�d���b�~���
����(���`�w<�c7���1���rbFef<��dI��>���`�0	�H5x���ݾ[ 8�n����d�^&�X�r[x���}�(���]Ύ*��ׄ�4�1�Y�����{�">>Q��(�g
�oo���۵���ԎaNBm��Z�Ȟ�jiJ�Z+U�Ch��k�V���B����*��Ϸof]�h���h�sz�E��L�2��xu��/6�r U��@2�ߍ:����@�u���=TQ�D}��G�D�6��M":#$��8�a�����w�*�T���ᵍ�fB3"s�p�Zx4���1#��U�a�$l��zE�[�Q��^�ߒ�[��!JP�(�J��Ak<���B�j����L��W9*D�Ǡ4�z����t����.�{���C8F���F�O_��T@�o�5���3a�5�v�P͜�n��LD,
tO.��)B��݇&ςz�L�Q\yO��	�[e��-�6Õ��>���,���A��V���&B�N7�ų,�7C��
Mx܎�m_��x�r��'�7 �bա�;�`�@E�J��+u���I���Z%K��e�
&5��)�K���}/_t���׫� =���d<�x=R(]1ˈR�ұ�_n��2d5ȹ��n5ׯ~B���[����N�W-�֩�X/G[m
����y��[
6��EV��QR51��hv��!����s��E�g(�x&4Mb�O�*�,��Y#�#lE%�>SƐ@1i:k��U���T�WT}����J�����}♌Az˥����h&�A������*5���Q;�˝�����ϜHj��iZc4c��+�W֣t�?XL<�k>�ȶ.k^&�0�O?�x�\���.'��ZLZ$�AF�\<���yxG@L�����.�S������=�f�[Ջ�W��尓��?Ws���q_$�F�څz�S�4zR�#X��+鰕[������m4�Qg&��w��6�b�;�B���̼s��_��Zm�R�]�1a�϶���v�V�h�
�o3D�6D[��:��鬶�N�c���u�Y��q�V��mh$�qB�S�����'��5��Ѱw�j�p��%�o��J�l�zY��\�)p(�������7y#Ċ�)?e��>��Ms��(��|3[8UU���/�S���&��y�p<&�r��eU�3��\�����n��*V6%6`�����1�EU�X� [�њ����0�;�{�_y"���Rd��L4ĥ�ܟ�vi5���d�X˄���;�g�m΄Q/g"�p_ʎb�����Q�5���3>��/K�Z+�8%���%�RC䰋����z�R,u�V���
n�Ow���%Q��u}�0��^�1������G�#�a��~��J��PY D�������x�s��8����V�|�Nje�D�X��Ʈg�䓝l"Q�+
��bW�_�T����u��{��TfR�,?��@ݞs�}��Bn�UVo�T�`?)�s�~��&E�7����>��/eR��cwsYѦ�`J��G��/C���g�j��!8v`7i	�a4�i��,���(/�̗�����+x���I��k0�k��'�8
��"�,�e�U1G������+Wcg�ޯ�- !R��C �]�gi�%R[c����zBz��m{*���FP�#��(��/z�?�äG4��"��v�Q�n��9[ٷ[In6���[���2_�O)	�I�gg>��U�`�Ӹp��`��Ʒ���k�!�F{�pN���Z�r �	���U�d�x�\����9���xm�/�:��M����XdAԑ�ey1K#��	�z1�rp$Xv��xՀ��"ОX_�imԢ6{���m���f��@xʓ\@��+�B�*�/	�Ne����T�����<L�K�.�F��`]�P�N�� k;,�Δ.��ENR=im�nL���{$���<:��݁tqB��kt�P�F�z���p��lKyw|B�/�#���Ж��&=˱ h�a�穞�HfE���|�G�8�����z�*�)�<r8��.ϲtd�W��*����Ξ��2E.��fT���9���
��j�.Z���d��b�1���/�@Q��Z̍���S���'�yxЅlc��젥	��0:Zڤ���%�6C�⑛�k��J�QIe�uW�i6٩

Q�|孟rM��[�Um5��:}X헼 v�K-U%hxAa��8VW6.�5����V����U5��˺Aȹ��JG�����~Oug��CS�m/k^�BH�p��a�0t���x�S|<�
:>���+��v���z̊��x�����k�M�Jx3k��B�s��D?֌JI�fZ�Uހ�$PU�m��54=.��-���h�Wb�nR�����FĂn���B�5hz���T��I�(�r������O��w>�~�l?�Q��P�2�������Cѡ�Ñpsw�S(a�H}��li��մ����� js~�Y�B�����d_�IV��wPT=�$���ם��@^M]��a�r�7_`�%8������U]�	=tg������.�t��ڱ�%����Y�xS�;j AU���q)��]����=���h�>�[�B���Q�"��wByF������-\v�@^�x˗��Z���dO)X��H�۞�D���s���:� ����[�GW� 1<	P�9�-��������2�>�l�c}�2f��(��S~�1�+q��|�����)"+��a�bm�̡�y��F�#�b��������&"�Йу	gB���X1i\�Rt�)W	�� (fK21^�X|�5�ʟ ��uO��4-8�^U'��(�V-��"�_4���.L���\t9-�愻������d`Y�/����9�	f�nq�cpR)��0$^X朙I�p��ė�`!
�`PF~a����t�/�7IH>Q�ȋN㡿=������+@�O��F]f��pt��ja��O��Ԛ���|�!�����d�q�L+���s$#�X��eI�+5-0���N�qy{#��*0H�#@�!�1/ǃ9�]���ͦ4�d_�L�f:�����$@�5�J��C�Gf�l�3JXPV��� ��I
����Q�Mߴ`Ky��䢁"�[S4���Å��!Gp�3cZ0���T��x�z�P�C�l��;#JJ�l�ѤJ�*�v܊�_��*R ���4��hY�l�)�0S����� ]/�����K�"�?r��Z�$�'�i���6�uz2v�[(1�N�)l�)������m�@�y�j�D?�L����՝Ck��3��X(�c����WGm����V���D�"$�_J�|zn�G���[��#�-��ed"��]���^Xާ�Ҿͣv� �Fi�!=i� �8����
|�xh!0#j!E�<�����=)o���斶����μ�(}��w,y��q!k���0�o�53��q�r_������/�BG�H5����0	�V�Yb����/i�H��{ƫ�7=P'�#D�q���R����*�3�����HHR�ڂ��NNa�O�Ԇ��� ��5T��(������E��W��]34���l�S�wj��,���u�q������b�N��SU5y!��?w����S$�:�����{z�q��Zű<�8�'�?�_	��8�0R��ũ�LH����<��'�X�i��&5���P��b���0���pB�JLOƇ�\��;SV�Ӎ-�e,~Z�f16�eK��f���_�Zs��\譱:f>�����y#̛��j�c\����,�Ao~!���y&9���Ŕ;捔y��>p�S
���K������qF$I��Ě�}b c*#F���?�o�2��`��Ph������#�A���m#,WW�QN/.J�>@��[��Q��H)j���֛ 2r�[��U^ν�>|��q{s�k�5�^���V��Gp�<���>|,�­.��sVI��џ�<:��K��S�dw^<�Ol�ꦡ��IP"�+�-�G�,�����]/�S�� H��	��8��+�i��uQy��3��:fk�K~46܍��tE�3��k��?\Æku-b��<�3!j�Re><�4�����L�O�A0��ݴ�$:�-,:�%!���}��b�{#�\l���}�_�xT�Y˅��{�L��#i�CR�61����=e�}����#6�=X;oOoA!z�|�2��/x�4��B�QB���"
��j�>O�r���8�l4W������sl��	:ĸ] �Hx�P3��*��Q�ǐk^-�S�\?�!��,��N���J�;�ZҎ0�I��GY��̈rp���~�ۤ)�� V�4/Ե��'Q{KBB֢|-7��u� C�S���r#�vr�A���(��VϱI����j�]"3�`{��y�{�.����1jv��oX�Z�V��;g��9`��2�ao#�6�7h�ǖ�)#�l�p
$a��v��Wn�iNf{�i��7in���n�F#��w�
5}N�y�4~)x
�p0��[Cak�6�4ĥ��{�B������T\��μ�!G]V�m�V�p��e� |��"�_��0(^2��ٚWꁢ��Uf�e�q��;8ILZ|2��b���N�5�/?���̰�'��J�;wZ5��0��� S�����h������ל�h�%a\4'I�e�"�w�>)��5$�\��4�d�*v쎫�or^]�
�/�	W�Oe/�qA2�fz�~
���(暈JCu�/iFY�c����$�WR�D<�5���@�L���0����e�܁8� _˟_�2J{nG��]���o���h 㖼l��/S������̎��Q��@��=c⃿�8r�%���H�r�G�
�V�,c疛�"�Fc�ܫm'�>��$�qk���>5�"Nw���
��6�s�qt�J0'�˱��C]u?N�eIB
�$�3zw��He�ȝ��^�j1���X���"2�]?>��;˜�Rv|ҹے����놅p�����{�kd���[|�B��>3�����X���l����N�7�	>U}o� D� ���m]jk�{PV�A:���}׶u�Zv�#!�`��A�P�] k��3���d��[L��T�y|;��f��go�s'�U���{�س9vz@Pv%xt���dG�Y��E��|�ý��9�C{LӁ`4�W9��+1�!�9 7��"ƦWۇ���,p��.r�[ZN6@!*hH��d������ݢ����iO���6�S��e��u����r|A��9貫m?�l����,�X:9�f�����b��а7�$�R���]C݂V��P��W�ּ2�_-�_V.���&�;LzҲ�HT	ʨ;�d(Ծ3F�~Y��+�A��y`t���a����E��Z��z7�_{Y<*+�;�3��i��~�H,î���p�'ۋJ�
�Z�ن����Qn\��J= m�*��P��/Z��é���Ե��>���D��a
(��,�����xNV���c�����ǵ��G͈�oo�O�-q-���#%'π�s���`Y���C�s�e�~'�n��/Ε\����ߊ�}�U�5�f�y�6�4� ����J$������˂�!}~�n��r�x�|uQ����H?&�h��=�=A�����#��F��Fr��B�Z�F��R|�)�X�9��$܉`q��ϋ�WԢ'B�� <�=�m��dn��_jV�-5�c������=G;,ڍ�d�K��#ZŐ��̼|�<%}U�<iq@��%����MB�ǈ<mmH���'�����u�媛�VKBz&�zM�K��v�|2�{iI��yN��\�ʼ�>���X���X�%���8 �|@���7���������]����s���_��#."��9��P4�4�#���iB�%�L4�@8ئ�s�+����T�=�a����O�.r��K��104G-�����)���q�jaZ�[<�+���fC���.�(n�j�mr�?.�t��Z���3H�<�P��I1������b�vXMG�~���������f$����Z�هM��Z�Rۮ��rT����J#q�;�`7|IK!��ȱ[F�� �_x�/꺍��!�X�]N*TX��ǫduW�)�<�
d&�*ӥ/˒�Ȟ�y�����މ���Mr+fh��w�}�KN� 
<#�]��:�<���!B�c��M ��-�V?���h8�͍�k���ێ�b�n��9WU3�.g<��)��%� ���J�ts�iS��Xo����d������,t�Լ`π�X��}_�X4s�9��f��yz��
O\#)w��[TǴF+I��ux)7w"��D�=�]9R�Հ`�u�?O�����q��G��S;j	�D�>f|:;�5���i���n+��mHg�^2�v��;������	ф�*��օ?��JQhlo84�0�( ��Ϝ��\\�a���XA[-�N�^��6D>��m�]-]�i@�AI��T���&pC�f�.0näF2��8����=�mZ�!��r�oS�u�$Y|��r³�<�ܶ�N�|��
ݰ�-��t�e!��C*���5#T�r�2ϕa���T&l�Yl8*��N�%�=�K�Db��ny���=�.p�88��-9U��a����د��7��v��R
��/
ĎH��5�Lë�MKÃ}��se�	>M����|��g5���� (n y[�EA��)
��i�����6w����3����,T#<��b٧ق���cDIQ�[���62�O�AE��w��W������'�Jqi��z�F,��Vz��5-jc ��~��Xwa�E
�ӹ����=܈N�%js�{�f�jl�p�E��$��d��� ��.*4�1sv�����D�ABI��[����J�ldF�1�+��v-"��ĳ�9�a����TA�uJ���HuX�M>[q|�eD�����5��%a��On�apO�'�r;Q�RLF݆� `��arm�V�gyS��"�ϏQ�gb��_����y�$�g="HE4v5G-����JGbW�)�~l�W��<*�\e*'#*���w��ˣ$����8q������M}����@�; �T��d�ŋ�[�柶]niNUט�6.=}��f��z6��iaD"�B��8����$!�Onn��RX��Z�(J,�=�:�/�ϠA�/Ф��>nZd���G�d=�4���WI�I'?�WJ�o�6�X��)�0���ů�Xc ��ZfXs�����?V%����ԷD#v�E6p��s����P:?�J=cD s
��ƅ����	Ą+�R/�k��c��D�T�b�y|�y1�*��Z�����AbF�͕����{+r,�B;�ӯ���P���bF��ڴ�V2�P4�;�0�丌Q����끖�2>$?�����c���)p��������ٓ_?�}<�ߐ�<�N��Ts�ܔA	�r�1�e��6���Bz���-��^�YΛ�x�p�F�z�$��.����]"��ΕX�K��F�߽yz�N�38a�F5���o^�.ߧ/�5�,-S���=�B�.�jR��Cr��VCYy��#Y~�7��A��q�H�6�0�F~��(�������d�侟�0�\M�:���&��1���V?yx��*�t0�<�,9�XGD��E�W�����3*ڇ\V�!����3�?f���m*�a�&byi�*�m^>�:� ʇ�R��g�O�'zq|��){�����/)3�޽y�}�7��B��Y>w�\���6�4bb�3��7��u<\�p���$��w��@!��3���<y��$+mXu#������Dj;s�G�=�`�rb��MȲ�3OW��FF�9X`f��r_��T��Qw���]�)`��Ϟ�TA�B�0�C��V�ǵ��*�/Wx��3�?�ܛ��Tw�ޕic���h�L&�i�%b�LO�K)k���&�d�b��o��]1g��Q�ɛP��j>�D�ʦ�F~�Ю����Rgh�� Q�cXd�1YtKz�:YD���ףG�6�$6@-�F��SV�q�[p�61�=������'��Bj$�C���_��qIB�Zݼ0�}�n�H
k���0�'4Q86�ZL�B�Ϲ_ 
2�K_�Ee��}[�����bW��� a8.���C�X�����%�Ϥ�~Qt����+7E���(���j۪M|h)j��JzӶ��X�3�Z�bt$�nzπ�ga�S�F\Ь%OwP)���a�Bɒ�E�D��֫Xo�b��Xw��+��ʎ���sQL]Y�"V��K�\#D^�K�kTzC�eحEݖ�b1�������#�����Ÿ�J�X~�:�I����Xs��jV�q�v@���9AIcW}q���F�9�g6䃭{�'�\{�h�Zn�4=�f���Z�rZ�`�d�m>�о��K+�ġq��q���/�ճ�%e��M��1r2B��I�0y�E�!���mR*#��V9�?6:cI~��o���Fĝ���b^��.���b�o>T{noK3ߋ��� �2� �Hv!>2�pdy܇W�<�M��*(�&_�
�ǖE|�<����h-�H���ؠN����M﮾js �Xf:����]���@�dR5�����WV>�2���1Vó�W"z��B�͠)�$���҆q���lՀ	B�����7pc����/qC�N L���,��M�����ĵ�ݍ�*BJ�%Q�1/�e�� �N���_�K��K������6�-���b�����(S;��o샠W������P8�����)T4�I^c�}�Z��^��	}Yk��lj�(�Z�;4�"�^��!��8[?�,
�"q�����^_��.w������� %}÷mW6L���f7�OD)Ω��[�</;W^�Vx���w~Lx9�?N��c���$�/fv����A�fx�%	Z��3)�������]�5���"��b]ö��4���YLp�V)+�&��{%O���;��4�+KvI�������>�ka��ݘJьRv���&0(��-^���9�o^����㑧���0	�N{L���!�(P��3���'/)jǯ#S�?h2k� �ܼ� �;��e;W�LH�MfHW�0����7Y�	r��l��|4�za�P��jQ�g ����UtY.��9k��>�1	����{��dx(�ϖ�y>��Z�/����}Lx-�ě�����b�ǖ�D���j��G�̲U�����B�.��\��y��.!!�I�H$ʻ���|}��qU��oF�/�?�ruo�`�'�J���=�>uF5\g���>����������A̪`5���Z=�o���W�
��\�'�?-��b��)�Q���{=����<�l����.��ܣ�
>�s���s�U3��Ɨ���L��睮~.���5��d��{�5�����@�:�՚��˗g8K2�]���]����[����N�*�h��~������>��$�݌Q,M矦Xp`�/vxZ�+Z��E���{#�!�t��.��;��x/�����.��U���ti��᾿XN��A�ɪ�Gv��g�%K������s2�U�>80V�����E��a��P
3�%}�"=
<�Z�n�p=L"�ja��N� �ج��dDk�Ef��G���0���M�l�N�C��&�=_�����&BO:�MS'���Cw����ʆ���u�!�c�����CAd�Fᬻ:���l��K��\��A�]�SĨ�[��Ť�_B>e�Fq���2�_�b�i�io�)+�m.�:�}F%�����I󭠤u4��A�Z ��ޖNZG.�mv<����;8�I�莻�pv�Q�?����%aI�!=|�d�����?�Bj�l���D�7�wlA���uP�Ms-$�ѐRu^Kڼ*��c#�|��!�9��rp7��o�������.�|����!%u_�2�T�{,u%Dv�g��)�.xą�Ї�e�o�j4�
e��ᣈb!5�}�A�J�&T��l��C�_G���I���?�TÎ��~��G�Fw�Li�Mz�D=�I�b��\�ц��T ��l%�O�p��r]�_�<u.W���3�!��T O�I�Z����a�dG��Ag�t����0woBL=�K��3���֪=���!U3i�]����#D��2j�K��o�?c"x���P$5�k���F�\��r�x	|t�o����������Lg�4��{ɑ'	C4TՆЁgM��߃�^l9�僔����_��r�b��Gv��ש�0���$��Z&�7���`��iO>	>_���}bb�c�~W���3MDx�pՏ��1��s+�xdI�.^� yL�]JO��iO}�f�����4������K��t;��) �Dj���E_N����c4�Қ��3@y��;@K�O�q�Kb4���ԑ����,��3	��wf�]l�'���S�/ŏ���FS�`��"A�7�0��ל��3��h��l.���!/5	�_B	��_|p��O�Z�)��ɒ�x)�����Q�S3ߢ��+ݧ��ً���gL|7LS�����m�j�٫�$|�����L�%��O+c/�o�^@ ��)i]Tn"!�l1޼����U�}�L(9Z?s�.�����p?�k]�'ަ�D�2���f�Ɖ�|����G�2Xg������>�}��pҜF�\�/�sr�W���8�ɵ�������c��&�wN�|���,�ѻm0gar �PE�!��c�Kmur��5��/~M��~?7��`�w�fm�%/�2h�く��Q�9	Gt\�wB���,>s1R�~�����G����H����Db7����W�}>8��Gw��cJ�w��$�������M�=������XV���-��`�aj�}�_S��H3�8�HC&j	�X�I6��޹@BL���@�"��Ԙ��#�$qi}?��epybzWǺ��t���y�X��`%������%U�`�RK��k�qO[B=��-�{*I��k��#H`&���7������#�4)�ۜ�m�>�s�t��J�s6f�S�.>�G��0#DU��-@Ph�ۙ p��'|~�p���+��#x�ի�	�W�e�m/c�̞5�e�E�Jb��x�[���f�&�;X��@RV]O�dv��k�t3�NR~�%�0>�
��A�k���2��nҷ����Pv�b�&$=nyfj�T$��I���U� ���a�\(+��[u�D�8�4�z��ȍ�\��s~z^Ͽ�tyۧ�t���"�G̏�W�����a��,����I���ʬx->����T���"BB�g9~ⰤV��/r4�1�`g��X��������֝x܉à�n�Wg��qi����cl|�&��oU{~Z�J���4>�g���T�� n#��0�@M%��~p[�L��ɭ���a����򲄪*i�2� m�dT���{�PJ[�E`e�\{�Kq�3`b'�JQDN9ȘN����fG+�<�b4.:]*VE�Iz̑z�W�T�H�\J̰j [z�_[�`.M�����p�!q��Ț:��o��
v�������0@���S��ZK���S��"�EE@�P&Ƶ߮E��t��F��n`L-�v�ߴv��W����It�i����\��}���)E�յ��A������� �lD�)�"7���Y�a%7�`$�e��m�gܸ��30b��>a��ʆu<�(�ٚ��,/3����o�} 3��6H��-��C��鏙c�ycs������XgE��R�5B�r QC�LBTX�2<�E�(��U+��v��x������YF�UP��NS��b�q��?y0q������x��R�L��X���:�Źf����l�DsGbS^�m�hԁ���П��?�Aw���N�C�epF5 �4�zչ/�;%$)0�C�fϦ|O0��6*����IRCˆ=�gCL%��G%r^#���I�1��HӃ�/�.n
����������m@C��ٴ2��\	ߓ��񾬴������kW9�1@;�m_�Z����o�Y��[��P߸y�@��0�v�AA��Q���]���A����@��l��3q�;�u�e��n�l�z��6��ȉl,�I����	��:HQ�l~o{wp�+����+jhOhf��\Q���cK�z��s�͝OӮ��
��N��C=Ga�%`�2]lg�rd��[&��O��h����>8�sɰw��G�����L�$�	xcXA3 ��5 1�Ǯ1vu R�FXUQ�qpn�4�
���˪8�j_�9�)>�牸&$��Ų0����2jt�0�;���7��"�xi�����;�S$<9��ꯆ��4q�ޭ#q��N��_�aCvZ�>��� 4��m �D=�Ad��䝅�p��0!W�6dV��I�%;tvWaM�4�d��ة��
0ۀ�1�x*��ۤw�s��u���q�!��=��O)���bz���Qx	/�z�1����pސ=�㓴�;D���o���0�$�[����fQ!��wi�Zx��N�����8�����'�3�s	�Ⱥ�,�'W��oФ�ٗ��*zU�b$��6A ��,�E�d���s��S�A��iT�cE����۬�?�|Of��p~����X�cW�Ҙ�gw�CS�ĳ~m�#�	�UB{F� �G�P/T.^>f��r�(0R�F��֗�_OԼ����+���r��.^�l5�܋b��WE���~�� Ѿ�����������z��_���S�
Xܰi��R� �/� 0������[��_nb�Ѩ��nA�Vi�8�"\B�fÒ#5�����!�+JM�K�7���Z��S4c �}���7W�d��k�G�Z#�t{�b`��k߯���]/8�����Z�K� ��h�-T<�F��À�[:nt.SPS���}^5���/��g6�Nr��q�r �rx��Y�6�C�y����55K�V :�$�(*���?L>f ��_�%�%W�o 
��<�>��6bQLL�V��N8f�W�C3/?�����(W��A��b��_�m��p��ޞ6�y��(���-��
��}�.�R����Wb|p���y�V��E�O?ȝ���Y�����jE�s		��/�;�N<_j��$�K�����9��Y�Az`��:ӟ�w��Qy���ߣi��o9���1�M���RB\�x�A=�U/���}[K8L���?���ۏ�q<��-���8��ka���S�h(��O�?%���`�������r���HY�>��G����~�(B�&�=r�,�W_�z\úr�<�Ӗ
��T���9����=��Х'j��@|YO˶ۛ&�u��UŤ�@Y(e��W�O��+t�������v�!xkk"��GKױo�*�[X�s5 R�z�w�g�K9^�X�!�+�K��t�!<l6��REf�=�4�i1��(���D��wa�������̓��+�1�ރ�=_K-�u��5c�A�L�(Ś�`���,9��e���z}�0��?=���P��Q"Z#��!˼'���w��G�����4l��Z*�G����X����{5ݔn~�6[�DZ�I$�P���h:�^}<C]D@�i<�E��#��n���������ߒ�z�b��nG�gJT7創Zgw_�\�1j0�+a�z�",#��f�*��%�Q����?��_���
�06��Ϧ�'��j�A�)ùRd��"����F�y���0f����o�ݣJ5��M�' +�Z�"4�?�$KS8{\b�C� WJ�Slj�D��	r�r湆�G?�R�_8�A��[ۢ'"f\�P�g�v�;\ ?7O&�6��z��|�Y�Q<���|�"�M��k{
���,�����.2?@�J���Oj��t��aJ�QL��V�@<L(�����+!�����s�ÊЀ<�,{D(o��k�7Yn��:[�Dt�;�9�\�1۹ն,F�t ã��w����i�;&����PƋ��_I,�v��MR����wrm>F���9]��~�{L�:YE�K��[1��i��1�V`98@��)Q#�s�_���$>����h�s/X�}��,j:݂��)~�畔�����dsH�QG}�(��[�;dg]�2d�:�/\)H�.ґ�o~B�gE)c�q�e�~�� �#�w�F*#z�w��i��y�:D
�WS�,f�V�4���J�p�iE��j<��Ho{E�\(�o\_�[z���c1��?�w���Y����r �vDwy��v�&��ǧ��H��B?h��ZH�I��xg2�X��e�`�N��O唝je��m�'	�kB���K����?�.�v`�sƄ&��Z�n�۫��2b��ᢶ��<�@�{�����&�<���T��G��t�$bMc1U��2��i�=�[ܤԔ� �`3�g����c��2ɘ0�5����JM�����P�ls�-P�@�9T�]�}q+�7 �%�+���I�ҍpf��e=뽛O��=i������>
�ٕ����_����C�A���ғν����+(&+���X>j��0�P!�EᇩR�:o�M��Orr;0�U� u�R`_v�֔	q�)+R�]S��X�_js5�ߟ/�	������f�k&2������P��F��_������ 5��}?]��碽,���^79����O�'t��d�c7����UP�U��"�&�B4��q�yg��;-<pz
4R��w�"##0xx
/�H�t5���fK�j,S�}�zR�|��R!���^�=ٴ��a3*K����a��tDӗ֫��M�80�#yΰ��?�<NKQG'��u��
�k-�]�C�~Q$�V��M�J�d�H����I>�骳ܴ�t�Xt���ߛ^�kM��/Z������/퍌�9D����ზ�6��>H尌0ɗ�䵐�����>ǆ�Y�=u�v�^⥮󱲅��CA�Z��N�ᆆ���@F9-�ǃ'׊0�����՚�y�7h�������k/nB5��\UQ����c��o��U#��^/j�>�8�!����# �pme�b%�֮�v�"C�������_��j���:FE��y<j�;�K��I��+�5௠p(l�Av�w�LP���ܼ�P(�g˺�(�1��e"F�OإJ�x�N
^LB˴�˼�{!":	��l�[�?���>��ꅉ>A�)`�.a�|�)�OFw�5#A�cۅnԺ��������1��s�#x"n�������uȧcnE�1|��j��6hYd�]A9��v��lݣ���������,}���u6�_F��f�|�Ew/��o'�~����<ts�I��N��{S/�,��R�\|q�E-�k.��9����賸�N��C���T QGz7/�������3�4�'Z2�`�ao�<�"}���HF��oQY3c�@[�G�Сh��*��g#,���.�R��E�c���$�@�[���I��weg=l���ݬ\h���~�J58i���V����B���r
�K���X2P�&���f�r�U}r�Y{FR�C�Io�*����X�5׋l��gQ�/	�<�0�g\]����o�.�� R9P{�8��؃�X5�d:ucv�y_���-��-�?�f��޼�q�Ⱥz�^� �+���_޵e�>r�W��/A�����@��Z�!�ͅZ�\��
�ۓ�0&l�0f2V>�JH,�Q� %jK�v�I̯�z������˨q���T�a��^����)���f�tXOA":2����C\��C��n���2�#s�y)P_���Μ��6lv����/����rQϤ�R0K^!hk�xQs"�(��
y}M �L�:K	����Y3#�E6�Sgڟ���1W�LPy8^�RhͤW%ǥ�ծ�}���qU���b���&h�6�|N�]�O7�t�����-NFc����Ma	�.��E�}ۚe�!��vN�λ,D1]FgPn�"���7�T{�4m�rp]��T��+��dJ���x�'Goܕ  �Q�>��2�=�R��T����4\l��+��K|��޶/\o��f�ko� �|$>��$1��Tn{v�{%}���ꁃ3=e��5˷�ɍ@�w�1�&�~�-��� ]��������� ^��Ĕ`����ڭ&���g�M�q^��d���\�f²��YS�P}Wg`/�.�H�|�@�X�q[K��.��n�{��d�ܜ���q����!짲��2|���NYb��M?����]v�/�F�!ܖ����,��I���&����=g.d�u��'o���-��Jd2���7����Z�^yC;PrR(l��ml� yI)-WCW���sA�`)(�P��n�+��C�ސ�1xh�(B�	���E~�\��	nY[
����~H4ӟJ
FD�3�_;<j�z�U8+�ϥvW���Vɍ*W�[����(s(*q��=��?�l�䔤\�iܻ�P��6Y9ٱ���W�!o��t�P�%����E�9��)��p�2&,'��WD� (�V��#cM�enSj�<wc&��w���db��h�y�֢t���PL#�Jȇ�u3s�!��z,��T�u��}�/�t��ZNnۤ�+��X�3��l݁���0�k@1sq�i�i�I������&s�<OSHS�ec���R;�=`�^��!q���`<���8���l�h��A��q(���y�����'1i?�V��]r��0�{�Yd�$��[�ᆩ�e�E���� ���K���C���'m.=��R.j�H���U�Jtlb�$���+��+���`]�h{���Զ@H{�f��:����^5�]����L�L�i�>
�����.���s�|� ���IV�g;v�oG2QkT��GK�ٖ#m
2KN/N)I���$�0���m1��N-��j1^5R֜b+���SE���W����Bg�"�O�؋�y��G��5�s�������J\6���E�kI���w���t���:3�km�}��1J���?	N� +5�و�R+��OOآC���+�¹�'��
��b����ȉiKED��H�C�T��:"�\���Z�B=AH�BӍ��9��᭕��p�q����tMT��C��/$��a#��u��'�=�=��J;է/&[߰�B&E��kϋ������@<X�;��xa��O0	4��0?l..�c���G���Q�Wb��(����Vw#X�R���B ��K]�o�ú��zN����u�����vS�&b�Z�^7��z��?�a-��c:�%.hR�Xw����V������@�?���+�lh����V�V@���'��>~��_:8@`�ǀ�!��y.��(a��Zg֓z�3��ib�W��G�c=�.�Z�X4�ɲʘ�.��䘓�a�w�z�}	�=�'7��B��T�z֌_
���xĝ8śQs2���E�|^�[K����m����!f���O�r@��(?_���4@�pqU��"���>ʽ�Pg�v��'�E�"�I"�/���.��Q����3����jq/[;�:2ԕ�ה �u{�XKd�E�<HݽI�M
5\k�U��ERW�n!���0᷺������o
����d ��7���
�=x!�^5��h�ݬ*�ޫ3E�"�v��`%��Y1v�C@��+y��8l�g�ܜ�,�����2���;�y"��)t�Ķ�@�ͧW����:�9��W�M�	l04�`^U�T8_�g�H�ߣ�8�	����r��)�)%.v���aٷ��#��ت�~%'����P��)�B#�r�X��co��Z���C�sv_���١i�B�k\(�p�]�K�YZ�N
��t�&�E�]���a%P��~�J�A��ҿ���*�DX��bs:��}�Ϣ@#�j��FYWtfX�Э��/A����N�Z�K�M��Cu����E`{ű�9�ЎB������<��K��eh����i،;�	� �5���MT����&K%O�%�
�4奈ԗz�EB%<�S�����K�W�£��sIUg�8�Cm�XiE�!=y3�y[t���-���*B7L�qCb�|�G����7`1��y]��E|�ޖ����$lӈ=�{�_��>��bJ"k�XZV���:o��h�rVX��}��ӈCJs?ްw]�;H����x�L�luz�Rx���c�� ާ�>p[�/�0<�p[	C��=�X��I��{Cu�=.�7�\'��yTkwR*�����v��HW}��X�2�C`���Z���7�x8n��LPFC��"0��7B|��Z��w����� 6C�1��~:&t�k|�ka��~\į������0�������������>{��\ c(�J#�u��z�iV��`jf-����O%�@]1p;I�k�H&��V�����IGu���=.��Gf+,)'�4V��!8�1���\֒pfT�O�
��B���~S������@P� �UB�^���2B
�g#���?�]��� ��^77���E}釡���;"�[<n�M�DvW$�D�{�=�WI�Av2>dZ~3��Z1�b�ݪ,�¸�N���ʋ�>�<DO�|=�A�,=�MjKE��%��r	���tC#�$#v;e�e7��T-���W��Uf�\l�֞&"|��i����h��L<*ß)�q6���+Y��<,�bN8P��I��/�n�C��z�@P�&M���X	YT��Xj���M(ݫ?0�s�v\���wݺ�k��^zV��a����O�U��"7�����lT�vo�&���uT�H5ΐ֛ '�F3��ˉ��~��6mTv��J��l�b���B���� 0�:��E�$?w�[��l:�@A&6Md��!mJo�*}�����b2��:����lO=�=NV9�yJ^el�т@���)�&���1�{��$��,�a�Ձ'05h��������.fQi�G:ip_Y�(9	UWR�@C
��H�E����V��{-�����P�29z���k����Cb�P�%����2�R�P�1W���Q3GI&��<U�1�tQ\4��}C�}@�ٮS���OTE�Z�Cg�9b[5!������w_{�%�g�cI�<M=�.��WT��*�м^c����j2��[�A0�mz%���+�^Ձ��4���^O��5@W���e������c��IO{�+m�q�����(�XA�x��Uv���dc#�u��]�X
�ԀP>_P: [:�����Xx����X�j���4U;$�^Ch�Z���*��k3��Ν�(ri+ -�;};rӡ�3��$��Z)��N_(�s :��D\��{O�T���
���%�*��P(F.�й�"Kб����`�����_��I9 �J[7g��=�4E<���?4Ng���v�����"uF=��>��Û�.F=���ɩR`ςc�D���}� �'�$�5�;b9�1�b��Y�!�8/��[J!/O#Ǯa�B�ik �Z&�B�������*&SC�A�`ժRc�'�1�`��uF��<��l����+p��ؼ[��_Y �������Q5�f6}hoF�xC�^�$�8����x�/Ը��U�n>wf��CF���E�v�l�s�cMI�y\ؔ����:&� L��D��˄Kdey/N�4j�[cb�W���8,t@T�JBF2/�53��3�����j+�6b��õ숱)���F�K ض�d�Y_�T��M��kr�i�S���C�m���	��Pr����{Y]b��q�2��c
�!(�����b1lb� %�ڱ�<�8V�$���8�=|n��/:G~4瘦���2D�o^2s�s�]n�1.Z+5���'��N�T~䨭pMrJ>�����$N�Z�C�<��������-�,KsX.g˃#>/cܹ#�fqP���H�Vgo��*D��Vo��D�с�M���v��=캦��<�+7#xM˼9��K6���l�Ŧ[�n ���Y�����\��������ǱV�<����H����!�ZBm2Yvr��/DI1�,c�6Qy�U���4"��(�lapC1�� @��'+�oMS�-Rm~�yrDs����u�'% 	ϗ,���[0����|Mv>�=O���ؽ���vB�$�5�P�r��@�_ �p�`��k�V7��"1#��kA��jE1���T�������:��i��r���kZ���d?��y�a�^�Oq}z5�2[�)hK��\(`��d�v,�h����~��{��Y�w+6,��h��p����]C��T1|�'�;n�7+��ܸк��U[`���gI4�w��✳���Teo�����7�}� \?�W��o���|,���I�%�B��;l+`(�R;�J�
�S3͞��n%*Eтk������w�tA<��t{OV�iT�O���?y+Yw��.
�7c����*�n3;��m4S�qUSK(�t�ʔ�B�;���3@6��ƒW�l��e=�MH���'��l�]��>S�B�gmZ�FkB��x���Z��P������X�{���}��K����ˣ�5�fX�O��A)Ln�L 7�k��p����1�P��^ҁߑ�y�����m$T:��C~�1�#5-b��UT�`�)i������?��,��êĦ�1��yw]�j�5�f���N`t
�~��'�C��tq�(ay"��6t.d�J9 �kf��*����W�LS����߽�#U{����c�~���ǦP\����i��+Su+�:���I"O����k��uWw[w(���Jy�3sO�LV���b����1�;Σ�y, �]�$)�����V\s0?��Ծ�W��. E8Q�tO���kc�������l�Rgsbz�>��ǿ�z��?9SX;����1�:0�x ���� v����.,Ӱ��.�yǚȺ��"*$3xNR7jE\r�
hu�����d��XU��6D�]��(���g��Th�;Ƿ,'��	�$\�64��Jd�1E�������ݟ��<&D�O0�ΦX�"IY �'�%�S�'�"&>�` ��2�v���W#t����,�!�ۥ�`yg�O<\�L�,��t0oʍ�F-�{Ã�1~��=���^!�m��(tr�b^��ǯ?z[�,w�ј͸�^�cV��?��{u�� �_��WraNX�rO,�u�(�L� � �[�_��:m�y���*�T��X;�M�}/"�����~�1m]5G�����HF=8�+�D�/-����l�v�0���x���Iw��o ޏ��cI�lls1�s������!��Ѳ�'��q
X쇈K�_�����fk�pȖ[��Y�J �&_h�?Cf/͚%��wn׿�X�^	e�z���� [�f�W�,��ό�AA�����Ep������u(̗��p'���y.���̗��o��do�W�+��g���g�E"wƢ>1����ԽU��qY������&�kgz!�e�ƚ�
mns�zŲ�"�gk�F������0�*'a̭�9�����+��~��Ơ5��۝�2�����bo ?�c��� ��K}�=�9�C����b���( T΅�D�ި�)�Zy���eN��B~̼�5%{�˸��;�.�7	g�	�S��	Xe���3p���|V�'\Ɍ$�&��U��/��IvE������
�𾏿xG�:����/�EN��`�&#AE\Į-�fd�2J��4+�T]Z+�������q7z	��0�{ocLog_��*����h���g����1���x
� &>�|Ҧ��KzɉQ5������ۖO⸮?�p�����0X�m�ii�C�<ps�n�Z*��ю#�+k�k�v��@�ij#�ҍp߉B��cA$/��	�8�&���'Yfi)c�^�^f}�췓!f����(�Z���� �����d��Sz��
��}N�1.N�S�&��<�]p%��Q�z/6I$��%4tp`�i|M8E�F�>
 ��-�j^
HYባY�ÿ�GE����wՠ(��}���wbjY�_�7�n=V!�Yݱ�iBѧ�� �RrɈ5k��%�̥���k�w���o��_`{-�Rr��=£6o������$@Zj���$@�-X�l^c������	I���֋+��D�	�������%�8�Ǜ{�C�	e�C�Q���|\|4E]բ�,t�ᛀ��5
h~�t^=C?7a�%W]���T\�PX��Ȗ������#�u��-؆��ܬ{�B����Wi�S*Ģ��w�~]m��.?��6�!�0�f�9���	�tVՁjds^��\�����,��z3�7���BR
�K ƓK�\d�̺2��Nǉ�Ϟ�ZiV�D�b���QNv#1�PO�Il��E��F���h�K�H��s��Fel}������o��7,
�4lu�v��O(� n����g�����[?�Q�2��A!�hG8�RF�S���>����h�d�x$���a�n)Fe���N����`�+D�㛆�R��~(V���{M��:�}��_(�]������7[�i�m�ҏl�쏰^��A}zK̦_k�:�hL/L��<EX��v�T`r�WA�p����Q��lo��g#�"=`���ÂF h@�/雕i����h�KZ��1��ω�.Ʀ)�cЬT=J7O�h�`y�j��ff��Ϯ%f�9%\�h:���~J�r��gs�i�<����<a�2��_AG9?�}�P"�q�iJ�W�|_�w�n$4$���Z�L�F�[\Q��FU����gkϥ�s�Z��ə�Ď�.�P����l5�uŲI���,�i�ݛ��c�����\���L9mZV �HiQ}�=��I�j��<��mW�W�(''�V���3�W�h�G�����e6��R:�7t�lv�/h4���Խ���A�+��,�F�����=�Ƣ7`<f>e���$nf�?q��9K��AKCMKW  �V�t��	
�U|@>�@0�� dY�L�m�1��n(4�1����P2�
e�6' kW��,��1	�5���IX(�j���jG��ۚ�x�VR�w���'�o����^g��my����C�t#�\0��X'aßG���ǘb{�i'�a��!@���m��@o����e��z�s��}V�c�.���;��	v�
�m-�v��(_c�ԲւF,\��`J8O�!"�����$i@1-e�r'�fӜ�_^ �fA#���x����7��t?بgOC��]1��D��K��cyt��I���b7:�c�I<�Fe���gx���s>� W��z�j���P���+ �>�u�V+���F�1!}|�4�ղH�_�<�*�J&}0�Z]��l��((R�����g�Aڢ��{;S�uiq%��W�-/Vw��i<B�#��
6d'Ҽ��/�3�C�ӻ��[�\BI�aN��z!v�4N��f�G@lc��#��\�����l��K�;��?��p��I���13Q�t�u�#�ʮ�B ���?	%��9-ܱ4U�o���t4��c����5�{�j=�O��L$���@��R�q���5�?�3������R\�	��wP� #1��������3I1rr�+����c=�>U��JI���u�23C;?
����p6��M����o������ӧh:뫦��bpʡ��PY0��Zո���{���5��5�4��&��#�c2��/2W���� +�(rFx��p�ϭfuk���ѭ��P���GoeXY c����˶���<��+DiZ���kf""?L��rh��A��G��y,jm�Ag�����E�m��<�~�5Nզ�g>2��	�,��"P�3)��\S�\Ol+��Z������k�1�i��OVE�E��@�d�%؎m O*�07/�5��~�f=J��|�?y_O�{|@��>Ap%
�#=ZG�%���R��CA,��2����c��j�����4����T'X��k�qA7��߸���g����n�d�����cs�g&���j��n��/H��>��{lll9�Mʟ	8��F�,���F���a��tw%�vw����U{L5hSᕼ�Fp	k࿖�v��	�tc�z#�K��03�>���/V#��D�o��.{�Kh�Z8�q�o]lV��7��':��L�sW����L��zY MeQ�c�4$�tĵ�1�$���R;�+h��Zfu�&�ܒrՇ4��@�״�	�ci˭��N+����\A�3�.�Q�4w���0�`QXډ���܋aj�Eye��A�7��3=����!���״���#?ǫ�.��O��v=��4�5�4�c�Y��-�eB�ب$�.����O>�,	�B�&{#��yI�����H��;�\Ug�2+I����k��e�,�^���H~oS. �m%�+�BY����-�x���i�i���/�Ge���M�\!ӝ_� �-$+\�Ҧ:R �᠂g��R.�b����V!����{��2+l�(\C,�m0��V�!�X�JQE͆YI԰�}��l�q`_ѩ���Z5�l���-�Z����h�,cQ��9�έ�I�E��x���S�F���κ|񀎩��ԥxK��>t}rpl�0=/AX��"#�ض��n.��J��WQ��_h������^��)��h�%��1dK �Rz�8�N(�7����Y��Z�yx�ǃ�m�	�v�!`1�yJ�ٓM���f{���*C��R���Wt�UO������g��d�>(���3dp��dq ����-�N�'�l�Ч�Ī��L[�Aq��|� �G(�����<#D�P���DA��s�G�t�L�UXd`�S��j�)�{��1���$M��~�D�t���A�_�/<؄�43]4E��w�^���|�Đ/���@-��L5�.���D�T���hP����g�^jkV�5$��Y10��F�6o�R��R�g/�H%O�"T��2�����K�Co:"��|k��QFJ"\5�}&g>'�6ӻ���N�a��,������h��G0_��a�o�y�|�[�,bG!��g3�!+��f$��\z�#g�'��8�d��[_��[����f��;�ؾ�_��q+d,������B�+����%Cc+Rt:�ˮ;璤�>د ֙�Mh�w�6�jnK[{dƊb$7Y�D�U�=(Ӝ4O$$;UZC���N��ޕ�t`A���=iy?�����C���
m b�~}ߐ��4Sl�wGy��ռ�/�@sj"/��Bx�b��d�<�OPYt��ض��IzzS���������T~��d�֪�W����	�"�֞�=�<���T�,w>t�|Ο����ş�a���E��4�p�w� ���a#V���+�����*S~̣�s��5����a2z���&����X�~$n�^H3�$�J��_ѓ�=�e�k��3���[� K�9&k�����߫g�铺-����T��O�%��p�}�~8��;��`w]4߄v�r4F����w_t]��r�޽��c%,�#��眾�OD�C��㰣�l�~[�3��`F��gZ�~I���|xp�UQ-��w���sȦ��Rz3?���w��Ř�<�.UA�x	#��ڪbH�)`�8ĉj/
U�|+@��ׂL��P7<8�e
�Q�jZ�na�W�#ɣ�7��������uQ�z?��� IM��;wM�y?��q���Է���1aF�k6�Z�h����/�cc�˃�#ejc~=��~��Lі�~È�l��yb�o>sݴ!*>�ĵ)�x 8y�ժy��������m��-;G9v���r���\�xA���q��E�߁� N���.�x2υu���X4�hY]��	�H�Հ83Ws:&���Pg��6ݲ�3�6��X���m��ǔ/�ޡ�/e���c�!N��L�։9�����O�P�l�-��U�j���
�������7s�E�7��w�8��`=�n�<�a"����HhO$��1Kf����b�q~�@	�$������)L�� �[9i�ݟ	����俠E���7wj,��U��S~[�t ��N;sV�ݑ�.j�p�YuqN��D�K���r���7[h.<�ξ������1��Dq�RL`�i���z[�\�d+�юI���G�#D;io�kWx5��Y �g�k�t�I!�Mi�T�{P���s�u>ߧ�.L2�H��/q:s9��x������A��g|�n9ãHUWP'&	}�z�'�'��i��9r6�� w��^�}>�s-MM�B_�SW��]}�=���e�x�������AnKp��L�"6Ɯa�Nq�53�����{96@+��|U�%���kf@�j�Ǆu��^��ލ��g��a.�o����X�Vuψ��>B���d�*��#��	�*�}�v�lp�=(�ISIC&�p$}��g�"�궕y.��;���	}#:����g�B�lh���ȵ�Z�b��>�Q[T�U��W!-�e�}ګǉ'E�i�#>[iw�ڢl���Z�꽴Xfk�����7��n��M�]����n^o<q��i��}=�U��6a]�3��mY�>|9��h����=�G��=nU�g��X��͓�~��njύu�Yhb�������(��e���:��~v��1?�ɨ9⭊��1AЅZ����
-��~{ߚcO�����g~Ҹj��ٖ�(������<��]s���q��&oO��ӏ�]>�������G�������S�l���f;���޿�i����<��ᾝl�}�~Z .p�9o٬�Nҁ��x�7����,�Sl��rn.G2�p8�̳�`.\|�\}�f�'�9�.�
�Ǭ�#޽�ǵ��!O���{~jJ�LşwG�.ˏ-�����Y+ytg��M����?KY��� ��|�j��[�z��Эܳ�`�άF��`G8/T����P���e1\+$֕)G	[q`�-_ٳ������5,x5�#�Պ9���2��d%�U�C|��ܐ
��6E�ήa�m}���O�\�PC�?���;أ`٨ 5�@j�����%��N�;���'�C��Bõ�j7߳�����*PT��c�4<�Ⱦ�u�O����}l>��Č��湋�����w���Ϊ}/�s��(&51g&a�b/��h���B&���Y'рG�ӓC0�y��D+;^ ��С^d��<��Gb,���:�prbl84r��^�_m1����MB�(���<N��;��:�{uڨo��L�*:Gi(��o�$������r�|:p������-?�Mmג�-\[�]|�
�A4k`������~���0�X *o���a�x�c�6~b���Kj�,�~&�f��j��WU���f�w�~�'~������׮�/,L���+��i!��g�M3��Cp�R���T�Ac��:9щ�-�g�:�?����[���ãc���͡~��սk��ʨ�vfP��Cg���E���6�"Z0���O�;L�@�/<�W��:����J��f`����b�.�I�	�-CS���R���oqU׶�Q�[ n�(7�G�B���?�Vw�ܧ%���Q02>�f,�A�lP�s'�d���x�㾄i�N�U~
A�F��e����x�Ы�=Щ8\Z���w@���2�|H�KS/UI�r�P=�+��vx�"�dBg�*�M�m7ӿ���-;��=9�E�	|X�G�H��,d�v���D��c(�UH��Ω��ɱ�˙���%��n�~���[�SQ�h��_(L⹉�Ϡ+Q�%�̻�qN��������t��� �´:��*
Q�?�g��Ry�8HS�g��';c�IC��948��Y!3*��%:���*:���y�^E�U�؊6T-�n��g]��j2�N����ل�#�C���>���D ��T�bČX"��pg�S��G`g��Y�4��*KQ�ױ
�����J��ju|��m����7�V�CB04�h��t�ǒ<��"A�Y�����.���"���x�Ãw�?���T�	)�ʝEi�f��[��EPHq�����p h+j��M�P�:R�\�b�!)��F�-!K�,Í�?����W���$~xm�t�e8S��mY��7�"!�
��FJ�X���:uM�<�:n���c����FN�u"��БI���k	���
5řg9�L�N��LSL�'���4t�_��\]�܇�Y^�a6�d5�2r� ��HsxΓ!�uNT��(�Y�jg�k.G�k�7�Ө�9�sR盜*�Dq�]�r羵b��W<�{���q�3Z��G�OqQ~E �Q�W*B}d�?������ǝR���K4YRϬL
W`|�mm���}�ͦ��U^��80��0SPE��dQ�D4�'>�������//���q`������{�؋s`��)�L��/�� �N���cX)K�x
��P�q�E�4�0�`;U�T�M�ld�弆�꣡&'�\����J��_���1:#E�y'#�B��3�[Ԇ4\L�7Ƕ��w������S>�Wu>��x̔7ǪY__�'z%�+��xױX���3�ـ>ן��8-=ۙ��;K|>�^>ۯ7+Ӗx���y��l:L���W�6��Y��_�=�N�L#x�'s�`��E�S���N%�҃;_���D��v"I܃�	��!�&c�r+-}�*�/kOY�ؤVԨ��"�}:�ۿu�)�[��H.L��3�C�A����s�bj�uK�/d���-F���L�1$��&��ur�FL�$�~���2���+��#JG��K�Y���ϲч��%.� ��=�B��%"���A�t�7R����#C��K3`:�㶄� ��Cq�1�s��xP��ǌ��'�wI��RY�I�G@
��ҵ���r;�7�[�M����{�|oA(5���ٰ���Hs1��{��,��)	4�TN�{�(tS�S��_:�T�sˍ4$0�Q��N-�*q4��\{J��:1>d])~�_ʰ�Lg��[����?��xCjbJ��xӿ�r��e�q�y��{�W�jS�l7:�CQq�P�v���n�*Ji8�y;(^ Z?�% /;����d��iqQ&T˚���\��U�C�g�]TQ�󷙽g8EYW9�7a����0�����s�f��*~�j�x�޺�\�L�3k!MJo���fh�n?}�C5�{�KH�C��$����8�2�����s�{��Ԑ?]x�|Tr�`�ڙ�{�"�Su���bھ���s�Ħ��luȺ7���p/Y���.��JY_E1���Z頑�[g�6,&����	���?��)�Uy_ #
l#���-�����m��4�����^���X��(�J�Y8�]��%�2�	/ɥ��b.�Q�H-T�Ç�����%H0�O�2�y�#�&�b�ua���-Cp�!\�j�����179+�����|���Hm�P�Ϋ�@��fQ�k�Z���R�aǊ�~���%�{y=�ֹ���u�Nk���yS(��H�y;�o�3��N��}�������9"/l�7�V	o�I�u+��V�F����tO�0�b�-�^30��_c�t�$m����4I �x1�uY⽪�\���bj���C:K-��L��a��[(e P8`o�^������G/�%�bЂh�D�ː�b*5��^��qh�j����u�����n�I��ڹݺƋ�DlΧ��n�L�b��k8�j� ,�/"��k����OF������6|�8qjw�u_�X���bR��xG D�hL��l��O����)�g�9��x��k(xs�k��C�j	��^�JR94�/��J�`���h3y�X��ٿ[6�l���8�� l^
�]F-��Q�:�q�r|�_i�C�[�V�,�/�e���z)�n�_�ƕ�߉>��qK����B:v��?�����rB���픸������4m��!�s�몐m�V��GL���.j6���U��-Zh�'�=29*6������iJ�2ψ8�-'��p
�J���Y���$���Lx+f���Y�*?\��v�\�Ɲ���B� 1�ç�Q�Vy���h>��H�|RT��0����*�kf���Q#��q�Y�i}K���]8������D�t;|�� �O}AϚ�[��H@�+����,�	ĆhJQ$k�f�	ʼ�~&撇�w�s����A��L��
� iY�rF���M��%��_z.#z�j8�'S)�TҲ�wcm�VoPp���e��f���N��'�*.����M��qwu67�M�vx;}=�U햎�DMɝ�]���T���:���m�]P�h��敏~��T�6р�8�z1�B�I��A����s��ZXH�`�<���w{� ������IKĦt��߹٬Q���!�T&Ic�,8:ǹv�㵽����`�"�9/��9�����Xo\�l��L���Nz̏2�<dj@�X�F�=��{��������_��_�ƣ�Q+���pNC�a�����3Dx�S�� ���`\n/i�ۃ>#���֑0���ϱ�2g�Yî��YAT��efi����T �Nm=XII���z=�{����v�k_U�Xb�L�_CL���*z�;�T �I';�
����:�c?�1�9��XD�5�7
���ՔD~jDi�K7�1�SBf��'�Z�K�:.Ӄ޴'+�N�t
�9Y�!��������s����,Y��E���g��Y�~�����F��-����w�Rf,j��U��P#ߦ_�u��|&�ηE7����|gS1�^����%А�m�,��і�V�Hq�H�m�3��d��XOR��׶��2��˳�
��Uc7k�ai?����Jk�!:�N]/�Z,����P*1�C��ƻL�;	�8�/u��k%�'"�w=[��z&�U��{�v%��K�¼$L#!�|�
�>՞4<�������*�s��3xow����ֹ�������+�Y!��Z�E09���"W���^J�J	9�E9�n�n+��8y��W)�:gY3�J�I+]���G�;Ԙ�	��`�L��죉_��m�0
]˘`������Eo&���aq��t�K|��x�g� 8�2��n��/�⑈Rw����V7�o^��X�qX�K�F���s��c�$��C�_�Z	�n�sMa�O֯峤޹x���b�q&fv9�i����~��P.�D6�u����ږ���ƛS��sTs�8l�D��)���r��z�.,��6U�Op�X�����Iv���b�Z��id�����AӦ�Z�����Q�LI�O�S�Y|�M���Q.���|��f;�����A�ߦ=+ފ�)�	V����\����N��B���ȷ�n0�zL�ς��ܑ��JX�[�g^B��{�Dܧ��`�|����ٷTޠ~�]$�^1�w��I?�]��{�F%��������������+'�0�.���_����c�,v[c$r�����E%��'�y\i�0�UK��|�&)JY�}ء�E� �'�WV�M|��kY*��	^���$��d�7֫P�w2L]x8��>���v7��#�IJ#e�z%�%\��]1���vz,��U�P(1N0���l�JRr<���	 )�C�.Y���9���P�A�*����c�B��4hXl^���D i���k�t���{6SMz�
BF�8Tl}O�j�D�f	t��~F!��(�.K��-b��L͗�M���	Oe?�pq���<��L5��[�f#\`-�DQ͟��l��H��1��5��G�b�E�z=�޷I��?~!|{/�=^N���F i�D|H����x �v����N�"�s�F'�w"!�Nz>;g22�A�}l���Z�?�GV��������/?y�W���6�-���W�c�1�<�RIv�J�/���ڽ��(0B$X��Ҟ��I���s���b�W�K�ꈖ�8����>P���1����3m�Աļ�7X8=C�\�6T��}@�5�	��Κ%~o�?��PojL�@�n8�l�Զ@�z��g�ɡ��~��;^K�g zb3��H<#��;����6�a�%a��tQ�Q\��iٟb3p�/�
��̟�%ɳ� �������C��*�*��R�<LPD3Y{o�O�L>����p�a��d�u7*#�<�"W��4����!�/d�6{`%D%�΢ZI�Dhn;�4�Z)<��:˒7�o�߭7k M�W��ULn��a!b�},�e��[;
��6d���9PчE����#��yPQ���Ɔ3�&X^�Q=��J����$�"�qHaǉn04T"tJ��z|䜶�N����G���B���U�q�O���?\�)��b��	!6ߵy���bv�=~��#	l�����k>�=����]�(��֒�����"2���XA���2AF^���G�/p�S�؆��y��*HQEbL&n�����.c������K�<���D_L�PA @5��HͲ��f���*���������n>�#��}>do�;���A���/����^%�x�C���+[2c#�4K��Bv����g%V�����
s���i��t��[ဇ!�W��r�B8]K���*�Dq���.��eq�4ނ�^J�h皐hwa� ��Whu֢�#>���P�?i��7u`���U��cp�~xms�L��'�\������i�m�D�k<�\����SK�#]���|�)^lZw���g4���R��5�9���TN&��4r݉�teG��{�QLy�j�j����/����ĉqA��,O���e+$'��[+��<B�݈�nS�<\��Z�����:��Ƅ��"��GM\u�������[��(�����=a��&�	X�'jS��8�ƴ���t. Ĉre�j�~�������&2Ě��w���ΙDջ�8��� �JǕ�l��kFec�9O���u�F�����"�0������ �=#g���g����$���gHL���*+S���^�_�jZ�����炦���pk#���좻��ea!��t��8;����
eS��2��vF ��5��Q����`�E�xo��2K2�W�X���H���'ހ�֧�q�&;Co��َ�����Q&�G�)���ׇm͊�
�#�F����A��O�Rjk��F^�E6�$�QQV����� O>�TϮ+b���vfu3X�T�&$�oM�Z�2
r�ͪ,�k4Ҙ�E�JZ�|�Hq�!�pt<X�w��i:�K�{�`��5��d=,9O�*��c��Nz����d�����'���oѶ4���[���M�<�Y�!!�������OZa!�#����qȻrc!$3�*���ۙ�-��#� m%���-H�(�����{���hM�#�U��@�~v���)�Ta�A��u*�IeU;BϮ�=�]'��YT�	D�AP"kB�#�o<6; ��+��1s�����ɯy�n��9�((2'R� (Z(��Ab�m�F��m��G`:����/%��9��.�l���L�3}����=�R	w�f4�8CZ��B�3Q��~w޵	�[�����üi1'�L�99o�g)whŰ���A����=�x��Mm_QZ�N���ݿ�Ή+��G�|E͞tx�T�T�	-\�?x�d
���:x�e�_?�Ñ�֧A��w��լ�Ǝ�,�9K���R�(��S f�B���ٗ��Zo����b�J�ǙxpP������f'e�K���(D/�g|P݄0t�^�G�.�����ff��ݳ��7*VZ��ީ(�z�~2/-@�<�xÉ�S��4%��^OLq�n�c��}�vY%�f�����h�Tb)`،�xi��O�FC�������&d����^.��?��b��y�p�����*�S�n���FZи��t���>in�:��*��o�p6i;�r�r��t�֗���f�#��w�U�0�3?��l��&Q���UY8�
WX�1�"�@��ʞ�����S�v�)}Nu�����w�r�O���Oa�J����4ݺ��r����:�D�ء�Wv-Ϋy�# �m �
�sI9.q�*��c����3��l�؊��
�-L���l��T�T˒x��|j���[������.�Y�'`mGA8��K�4����7�A�*��ֿ��S} LSmo	�:�k7W5��IS�-���|��#�;]�u����Ő��P��^O��t&���t"a�1ݩdm�'>�M���̏!,�m
���0��&��z�~x;j���|Iř�����<�6��V{�8kK#��*;�'8.'�����h��ʴ'�m���Զh@���?sN��,����ȭ^�c�#��("q�n=a�f����V�dp#��~��y:�����qR#��p���T�]6a�,e�����F��OY����-o��`"Ł�H�%.R����>�d��.��k�����J�����ѢοPTk�H�i�K��
�T��@�"����o<w�a�:��u���ه8o����}���X�n�oX�p��2�����K����f�z6y��|��<˒�-�Nw�[���_7����RL�|��V�����uzPBg��JK�*?�����;b�-�]K3g��:�.�U$����
��^	�B(f�!����^��%�4
̆�i�lkr�L�V�lc�����e�`n4ه��1��F�c���=�&瀿�����s�I���t��Z�-j]!�쇓C9Ї��t����1�\%ꨂ����I�[!:h�$�>��V��8�h	A�0��I0ޛ����d晐��5��u>�h��X@��}�(��~��
Q����U�\(�[��:���15C4�*E��0�q�R3������m*��pu�T�+�jS7�n(fc�����}Td�D���0x�:�Mq����l��P�J䉨�F����>���:ޏ�������}D)���2^��.�c �e�A�#N��{H;H�n^����m��x����������k�m�2#�� �
�҃���f|e�8�q�V���4�Y� �$d�m�'|��yE<>Y�'��W�(�'�2���Y���=��E>�K��縍X���	0QZ򄺡qf��H��wl"�]�\�ۜ�@�aj>hC���w��,���`0����.�p�9��D�,����%xV,k�����_"��Fue^���g�=�V�Β-8��e��\+�(3`��LU�Xm���< ��d����Wx�V�K ��n���a&�Ԁ_,e�jC���OI�0�_��]k��/	>?�D��+�A�ʣ�U2�2�&��<8~�;�܍�m`��JPe{�	�8��g�s��G#%�\��Z�lCW�ۻHJ/-O�I�폰���,����.3-���+!�I��F>��a�HRL1�!���:.�
Z�<�q��(f�'b�q�u<����!
��@2�Ip��h2��u�K�MT8�ʦ<7y0��b��w��Z,��K����qH�OAX��]E)�1ѸӪ�L0- -��%�O�������P�&�\0��3����o�j|Z��>����"
n�+6%�wv0�>�r��C$~���K+�����$��N�*��V����VV(# O�J�%��������e�y����^�znp�9��VST�[�����;T����D?��T�=+��D�T�]��%�u��#pJs	T����yۓ#�V����
D�3g�x<y���͙�>�Yj[��LW3�����Ͼ�����?�vN�W��!f�� �d3擹4�PT��;A�R���J1g���,���tG"Ʈn��і�ɽ$g��%�t<�pM��<�!u��멠�K��'�R\[��ji��r����K������=|��C<�v�m�;���A"�̶I��Ư]���+������v}��t%�_��pВR��!��#f��jDW����n�1�$j7��ў�#Zl���+_���ѻ�M˲J�jA�l��
ǾS�����_9�c�ʆ{O�9��J�#��|�;��ٟl|�,?�h6��`%R����ҙ����
�p�x;��,\#�h_ꡜ�7"�c�;�|9ø�tώJ���N������������uS"o7� J��b�� ljr��ŢI�a.e�m��;�ت�mYҌY���ɋi�p �_^QZ�t��TLkRY�q?�'��F�y!=�eY�S��������y��/���xǰ0^Y�4Y������d!����1`>r�Y?e�Q:�*�	(�/���i����τ��cm��������MQ�>�o�[�x��5;X���BK�]��)�W6��tԓ�jI��I��Iܰ�������E2��/���2�}��+pϮe�b�~����c�͸;�(E���Zg���Q�z�4��C���_l%��{��D� �S��o�M '	���xHˊI����G��;�r��� �+��{�B\[�h��tT}�MOFY�k�[,�zm(��L���i�x��y�;f����,W�R9ŏ˃����O=%m�,k7�־����X��0+�&;5��u5���nO(��~SJf�O�I�&=��(�r�P2GS"��f]�O�[��Ӭ��Ek����n)$���p���&آ"䊩�M�e_��D��)�.x��6d7�<���x�n�q��s�Z?�ٍb	�4gc�k�Q���S�ב�͹N��>���t�Mܕ���
��hO�bb"�� *V_:D �����q$��\B��A >+�p�r�5=�1��z���8s�Mʖbd7�Bg�$�.���i��̍�K��"����h���y�2��c_�J.��x\^M�6y!62�(ݗV�6��vy}�o��zf� % �V=��mYaAX�R��5�{�t����"��sd?�P���~�u����	���S��u̘,K4����D���U��$x^vR��7<�`T�ֈ�}kvV$��s�@�v=]^}#�n^�,��z�D�-�ȝ}OI8@�MO\v�\ΎkBn샶܄�~u�$D1������6G�e��|����p�J��CLCx��/���>P�t1��=l, �(�N��~O�,�9c3[����wM@Ou������p�R���i�C��$�
��:3�.���rt�K��5by��R �fA��ݯx����Ü�}�3������������?�{p�K�7��^���a�ڀ�#��>�-p?�L̻*�+�0��xT�N�u��w1�Nv����>jy#��>�K�<�ˍݧY������cD�Jy�A����߀��:�	��D��#2��t�j6�.�%2��Y�)�x�2�7�Z���fA�V��t��Iaж�
Q�_N׎0K��>R���R���6�8 �U()�+�>����ƌ�{F����XK �7�<tM�a��|˫]
�μdhR���>�l��λX!B�;�FB�g�n �b���B���P)xi��+2%�(|r�O���>�|w���rΫ�����$;��c_��&H3?ڮ��I��6OY���O��V���)P�@�Y>B�>�w�s�W���qC��٢���6��>X!+�:P�)��˜��� M
Ӎz��e�$A��-�5uG�g*˽���Vz|z�w���A=��1���+����s���a����9͹T����I��w��o�s�>r��D����;^_��^E+@�������4���[B:o�ko�w�r��A^,;�{O�b_�eu���0k�(��#m���Pg~��d=��
�%Lݦ�¥h:4�qL���.���sA�:�����Y��6��#�c�!��q��s`Z�g&MA�bcת��Y0}
�a�Y�X�ΪG��nj�D�T7���*q�̰0�F�Phɬ�����D���p���p'g�"~����9h{j���vX~_�^Q�P׳�<�a�l��װz��vTnGp��gjN���Z�0��KA �Ԙ��d�'����� ����Zc���y��W�@�Č #b��q��W�j3�$-��E�^H�s$tB]���^1]�9�������� m~�#l��b�::�l�z�z@ՄE���'��RV �F
S#�����Yo�H7��EHԺ�['y1��(�[7I�&�wr� �3r�I#be8�b�XH��^�����5��u��
Q�:9Q��Ho��m�� �/�M�-�e~�'η%�*�k��|��a���=�[	s����l2�k�J��i/d���4ˣ�zf�ɳ7�R�K�EGo�X�62UN%e��:���)[--�e.�u2��DZ�7A��&,;|MCQee�eq>�S�Ih����g���z&���3����6w)+������I�j�SZtvȎe6���V�N+��J�2�"�;D[nN^ٶ��8��#�o�{��3�d@��G�j����kA5��]a��6�q(#7'@bS�F�,bIu��rx�.�ۄ���6Zc�W���u�bӳs[�b;�9	�)���߾��Fnlֿ���U��Q���Gج�`v�
d�C�2!������d��"��pH�򲥉tݖ:�i��c��xc��S��nqm�B��,#��M�O�A���3\+����Z"*�$N������9��%"[�CZe�!eλ�x�%�r4˗�6���J{rl9���� ��t6h�0h!T>>�z��!WB-p�Xj���1Nt��k��F����kD��@Χ��0����uʩ��}xB��}O�35X�]�$>~Ĵdz� ��kmJT���D2���>��{п���	C1�&�߀'�7���s�ZՉ��XW����ށȆ�K��h�U�d{�lq�}������0av�V�\� �䷻k	�]��;��|��Y �vثf�׭G�-��鋦�b7�2���ck;=��[��`�f�;H�����R��NҐ�B�0�HC�q�1���f2��_.�V�c��;̈�>"���0� %&��CKk	͞�H���GZϔ��{�X�q��tۛ�l�S�?�5���An��8a[6E}���?>]Bؽ�*���j
���])1�
����]7KU��۸�{	��F��>wK�q�)V@�,y���'��^��BAG��V�&�/ �d��8kh|3�Bv�Զ0�ɧ��e�����Z"n�m����U���ɜ%��+M��)�C`��ϰY��ۤ
���@��8#�A��0��L����hcq�$����,�����<�XN�,���0�Pwp��u�~����Kȗ��Z'Z�����~�*�A��n[���.����K�G[(J�f��K��m/[aOS����d#�k�.���I���i�>`+�]o9xz�^k���^���t���������@��)l����i|���caIY���_��`�7������b\z3�u_',~�N_ɘ�,ӊ�E���Q����(��1wX��G2Z�Q61��jT9�aП�I�#������Uh����m��L�{���R���آ^�pP�Gjϰ����!�"����@J�fN�3�",�>rq�3|f���P����t$��'>�����]��L,w���-����9b��J�!~��>s(���,��π��ߞ�>i�<]��&�Gj�;����VA\�'9�0e�򗟨ۻ �f�	��K�IH�N��׉/�0X����7���k�6eu�6)[V����ѯWDg.ܷ3ɺ|�f]��sD��o�?�h��v���AK�	$:hɞ����M0����=	�K�D��,�3po�MȘ��T�����QJ��~�l�!�$��9���n��ݐ��@<�͙�s�D��0C�#"u.�9A���#���9,,���I/��<X�RQ;ؕ�a��d��<
dS��Bs�	�B���t����+)D��`~�8�>7�:�)Հ�!�h��� Qw�a�<���@կȰT�{0���2��8`.���f6�= F�:��-�A�q-@)Hf��sp��+�j6W嗓,�/q�c	VW�Wf݃-?��`Ԍ(��昙���P7/���^�tͥXN�J�D
]�1����KT�9��0�u��cdlp�^����d�K����x�ń+��!D�g����F������N:e��č!�V8�70�a��T��Dn7ŧB�W;M����j>��	��4��{�H(�1��>�����O���v��e�����z�
o��$_���E�a؇���'�z�'�oDE�bzwG���S�V]��Ά��P�dN��u�0��wV��݊L�Hʜy�����ll�h�4��@s��W��Sݽ�z��K���-< G}�DHa����v����)c����1�w�pv�U�x��{�[m�k��K��"����9�G��S��E�q�`%+\>c���x�.��	�f�R��-���%-,ރ*8G���".���i�� .p�56����Sǟ�eh����5Y/�Gz;���#�Y9� �����<[�bJ�ia���R���ꚰ�+�[@x,��T��M���'�t2t�,��L��d�5�`����D��Y`�����.�����ys�D�eBP�y��V���V�<M�Q��g�j}7������_h���&3�C�q�	�^��3SgQ��pR��ѼK�4��:�l�GN��뽇�ӷ���a]{o��)�(����~C�>�	�24P����׆k�3hӄ\�{���~V�����}�Q�գ���ny��}YПQA�%�#.�+���
ear�ms1���q����$>G�����/�bs�͵�����ã^�*^��3A"�������M׵��U��Rr�����L�m;�=T�����\�q��OX'�z���6����֠J��sp�jե�ڝ��$G8��^�	�u�j��Ǚ��l/<\R�z��#FE0������B�K�O`�&(���/�?�>E�j������W0B9�n�sL/5uo2��*���nхk;tts|���a�V?�\c�yR^1���y�}�>�\���Ńݽ�#T��(���%���U���@5!��(�i�8/�i��_"K����\M��6Nϙ���3 ��9�2T7Fό����{ᬠ������ ��ȣU�m�$@g��2	��2M���N�i����dΗ��S��� 2�,bk�J��)���7�;�N!L ;��Oq� 
��A�`���9����7����Q�1}VQ��_�	"\~x�@�Xg�c̿,����ǪM�	Ġ �Z�ߠ��B�˴�5����iۺ=���>]�R�<��
תf��Y�{�b�K��m�[ kk�B�+|I˜P��g�����W�#�ư��_>��U��o$��M�M�A+U1���􉡺����Hͼ�!�N�(�v�a�GK�Z^��#�&���Ȇ>V�}#:O��Z�n���z8Q�p!��Sݓ�W��4�S]Mѧ�d�Iu����)D�+_\�%��걘Wâs��>()��z�y�s`XF\��dfil��'(�+B[E# ��D������8Kn+8��Sd|���/���*�Q��M��/�r��]_jf;�z[�
�_T���U~YlU�J�ن�Kk�y38X=�W�� Bw��{�"���^̉���i�ײ{jQ[�{�g[�y��Y�qm�>-,Vْ	g� <)�D
�z�o��_2J���eQ�w����&Gw~Q�����q5��Vu���j�r�m:͵��lX���ܱ�v�����<gcP��'����P���㳨��ow�_y[LPRT3�/��~���lB�;�p��Օs&��w�}�p{,f�Q�1{.'B ?����{'�s����;�\��䯔���y��jۢ�R�M\������g��h����!�﷉4@��<�`�}+X��*�DV6�o��B��S��N!�Y�
V���*�o1k����y�Y�X�!�z3�e,b����u�!t6$�$6�&U�V��̌���aR�R��X���e������jc����X�g6�s�zH��w����<s�[�[�8fƫ���ɣN����5d$H�{�9�خ�5���� .-����ˋ! ��95��d�RY��Qύ���r+��h���ШM,�6��q�o��������ꇉM�;D���4�\���78,N&�}ՠ亳�q����i$xD7�o�wV42��vV���%W���{����E���r��D��v��v�Y�#���[f�DVP��̴p7����n��;!_�w�j�J��0�����:���F��ŗ�竰�����S���4�O����\S`/Xs9i�CF��*�It'mᨮ��w<�LΨ��@9N�N)���-���h�؎�3�x���TW��EL�.A���H�jW���:P��ɡ��!ϫ�MJ?�S!��sR��#|ϞkQ�W��E��}�ɑ���$2��Y!_�Y4X�~Y���N���A��WP�"ޢ(�m`�מxg����r�dH��u���$r�qu��-f"�J�A[�7��B^��  �!F'�[p�Nz��H��9�sNn�+pky�]�-.�+jxV�,������|��������� .��Y�Ϭ��������G0��
Cٓ6ȗ���lI�� ���9ե�2��J ��'�,<�F�o�O��X��8�FT���+�J��_i�m32��6�{	ކ=��Ō2	RV����*(�G�����L�G W���ƪ�������L�Bj?�k:�����Z�zQ�P<H�-�g��%�!>l(g��GH�Sl��h�vB��H�e�T��~�y�)��I�و'�oI� /�߽M��<
��̠�<Ln�1ēaeN���Ò, ^[U�d�r4�0�OF|b�$Q�����{�CC2��" 3����ҵ_�V��NAL�+m�5��.��/��+K�{�����a� l�Yw����3D�E���;�	�w��ݯ�< g��\ʙ��߻W��gb8?EU<���2�X\�C���Ɍ���g��'�t������M�����<j���6Br�,�mό{�L�j�#�bFߴE�oN�~�u21�|^2l��
�F�֕�p&�����B��FPiw�F� D��Yo�	����W�HHcn���B������q���e�S} �\��}�N�_b_�y��T����sĖ&Ӕľ�R��@�܂��(�Z
�%�1���!�;G�hX�t�8�55��e�w�:��M� ���ʕ���&�'��h|�����I/ ��������Ƈi^%�ȭnެ�Y�П�/6`��,ћ����a#���a^�>wpi��-F����<Ǽ��WkC[�H8�˞P��P�K#����p$�ޯ�1�ڐ`�uq�\���3��h�0j�;�q=�}�3Ip���{�K\�f��O��q��a�����no�e�:��Zâ�UC���TE��`h�UŌ�-x�D�w�MDwA_��������Wv�(�o�N���l?��SR��a+bA�p?e0���,��VEvgGn�P�bg���(?���;>�8AIF�U2W��)�&�!��{^��/����h/�"�d} ���&�Dm��&�x��t�h4s�%�;��+�V����T��4[u}my��,�Q��Y�T�d��W��sJ��%/��I>�Ts����x������:��!1�UA�[/�MN�Eu�<���N-��e�n�0��%@u�~p`$�-�>�}%1���6#�Hop<2�!�1��7������B� ���E�s�dR�v�4�"�i�ou��
�a�@-}�s�k��Lʣ__:�"����1Xu�+��=� ���<P��^�U,S����ô$(K$�:X��ɅJ����]!��
�Ӧzz;𙟩�A
�m���8!����z�b ޔ 2���1�O�{�ayq
*�HB�q��ލԜ�h���P�ӊ}�� t���y
W��o�dUZ�6��.ڑV��9�it���j� 6ܵ���n���W�n�Ɍ<)दYЪ�F=+_�%�bi픡���=k�zp��|�hw6�v&x�@!7�H9!���KR�{�
U�CJ�4k���f���uՌ�a�z���9C�G�1[�JϏa 0(������ͧif��A�����6�{�;�����U,[>H�����c����XH�az^ׂA=��͢5$����Z���wD���lEվ�� �D�՞�������mh�n���GEm�L�a��$�G��r� un7�BtvhR�*K�#Ղpm�%P����a3&)�54fS�za12��SŮ,�+���]�O��LqO�P/�Y�oV���{�1�^T�_vb蜔�#��,��]���G���?���A�d�a���m�YAf����!��U~������,�4�I�V�K�����n�/{#�f_��1{5H��H�D�ơ��")�ߞI[�!UK�x0�ё$��&I��	,Sф)���TY���e�aQɥӜX6�Q
^���v���WQ��F�5]$��DR�5>���zsv�X&fW�)�S2����04P
��Z�Yߴ!U�S���;�[�]}�޿y��Aw�Ʈ�I48U�i��{�N7y�|LB�`nY#�&��?Ȣ��1�������
5�4� �8U	QA�H3`;��(<��#�;Y-B����Ř����c~��[87�j]ֽQ�m1D��1ǯFԥ�JPC�������+G��4Aw�m�xG�w���3�P�La�s�V�� VȥL��`źq�{Gt�J�3!T,:=[���uVl���pSEw{u�pf &C.��L[��������I�H^��\�|L�*��i��hY�N��a!=��^~h��x��n6�aUL���Lz"Л��Σ���0�o�o �F�9�7�l�2�j����9���d������+����+�\����WJ�:K��NF �k�c�)2m!���3���u�R^�]������<^wz�D22���N�ŵjn\GJ[r�ò�7��.��j��U@�i�K��c��B�s���V�-�cD�����2�LGְ��^"�\��f[�r��0r�ȥZȗ���q�!�Ȕ8fi��7+Z%�����a���e�;˂��O޹�8 q�����p\��=z�҂��pyZ0����|'f��S­`�ŋ��DJw�t�������d(��V�^��`�Ù��D{?�}�lE�3A�qOQ��?��\e���+œ d8G\�Af4�| �e�l�hp�H�_�4bA�&�=������>uI��7�P,�<��}	/7�O��x�ֲ�V��}��D���Q��s������T�B�㣥D�顉�M��qڴ�^����p}��Q��#���l�p�~�ǖ4��.ԉ��!���-Q��s����a���6�[F�ad����g�h��G
�������Wg�	Jēn��L0�Q�hu:����]*<U���%}�����ť�,m��#�L�cF�p �_}*��9�纣K8�ʡ��.e0Q��oJ�+��� V�/9��]��nl�@�L�j�A��"�~N��g���{�])z��	���i��J���:M�:G�&T�i�������<���3n���hy��:�hĞ�S������p����}�1=�^��n���Q?+xBKݟ�Ϩ�搻7��]�����o����B�Ǥɩ��"�/c�ʠ�^.��_U,r��n�n�p&U���I&-M U�E��{o�(\��P������ik��u��:�����=o��판±8mH�$�.���G:�a�4ˇ�4IT���v}.���7��˘�1���;,L�Ֆ4#���jRx�����P��tu�>��C1�	<j���S_���G�s��p���v{�;��
>Y��(:e�I=ćKƬe���2��f�7�2��@u�X
��J<�|GzQD�=l�uΑ���y��E�b�,E���]$iPP��I���=�H�j�2<JPHҀ�
c���]ϋà�jm0��&pС���,`�4|�EDz����3�N6۷]u��U���{(�#�wDw��j�6�*-O/XDγ-Y���A�N��I[궬�����N����Q��y}��E���f��e��3��HA'c��6���R���b����O�_��&I��;P�@��q5k��G
�]8K��{��=�B���o%���<g�#,r��:�p�[ہ弜Cc�1zi����$��%h��6[�$MK�u"�XX`����{�\�n��Tk.�{����_6	D���]�W��%a��������]�Ʌȳ嬓��ȉ_�Lq4M�i:�s��V���a#���퓃%���y��xU�l����n�sم�5�����)d��h 5��z���'�G�135�FO���$RIZs��i�I���I�(�����6cR�[\B޸�{C$�D��fe�]o�C+\WU�	�OQ��-}�v#�1)��C�>ƥ�:���%a0
t�4���\�N%��bK6~�L ��_GW%_�����ػ��~����w����a��!M��`@�E�"��"I�T,�J�g���c;ڭ��!�MK5Ţ�T6b1���@���U��_nD�ʱ'�Ơ>�o�M��Ʃdֳ�'�񂕛"6z\�բK	�r�>'{$Z[hm4��v<~Ȝￆ�rP�%F5i�9�9�d�K�'�R؅B�dj��k����<�\s��8���O�IZ;��K��'w��{�(�A��q�,]ĸ��DD��c5�	�]�l;���ߏ�
�R?���W{DN���[Pt�Lo�N�,����,8�5'�β:"܁��]QF�c��3���t�bH(����������d��q�@�\���-�ŏ8�0_�#Z�A����d���T��6�W���Âa'2�c��*�nt�4<�o�S��`~=�����a(3����Z��AY�d���a�b�.�C�2>E���L�����M��{Kk�ϛ��ME��@l�V�I��e� B��]�6{w��q7R�XQY\؆�������q�A@�w5A�O\ 1�	��_�yw%�!�[�;p�G8l�aK]��LJP�(МSubZ�pV�;�\�wP��	����do'O�2�mL�,;�W�
~���!&8 ����qv�N �{�1��7�ø��B`�7�?��pą��M?N �yl<�A�pX�wZ�R ����� �;R�T��q��OǠ��s1#W�ʜ��j�7F�7��ۆ�	���B.�!��c>�UiD�?�R����m�UE�.\��Q�Vb��k�H�!������ ��Sw�O�	������O���Q«�j��~��/~��A266�ں��>�N���n� ����G7�Uƶs$O=��g[C`��*5�����#����2�f<I��}�k�!ݚ�P�<�>��Y����Y{-��E���O].��,�u�7)�<�mjvz�(��K��O\���䨈�H7�zi�-7�g�ľ��:�u
��:u%�n%�,呜Jh�`�����8E?&Jd�v���*��ڰ-���ށ���w���'�>�:�/���x��ٖ�;�19�2��X��J8�Tr.�c�N?lT!��%@����źw�t���=�� .�����p��5��)a�9�=�Ւh�[#�i��X����o��o�_�M6 2��
�{DECp��5L���*��j8�PFP?�T�;`A,3�돔w[d���N��0��l��W�4B�����	/���Ѵ>���}��%��G!�ߢV��=&{�
9��-/�A?)�G��0����hN�eò�?����K���T�&J�-���8��iœ�A�՞���+��w�aDG6<̮�=txΚ�����]"�tL�*G�uQ�^|Lީ�4�&�2� ?���8Շ����P[܉?{�I_� ��1���Is�+Z��Fc�E�1��:�!:�ħ�'�}�Cs��q�ܧ	'�W�� t�LZ�a�ƒ��:]�K���lG]�WX~��R�0&o��X���G�K	�o�h�� "��(�)��Z���j-n�?��$zYL�=�>��
�Ĺ���r���*�z���}�@1Jֹpgy�f���d(�[��(��5)��򒬕�G�1�}��6M!\�g`5����b(hl_�d���A�*�?Z72e�� ��-��j%ֳ@r�"k:1�d��Lo�D��.�|4��m�+9V+�P���Yg)���n��c���IR��O��9ڇ��z V|��YQ���d䘁L�C��A)J�e���7{�z`� }�_�(}�1�?���m�I�5���vJ��7�����m�����N���~���xpm��y���۪��%�.�o�g~�%�@�_u_aO����DW�C@�Q�Y�C+��!Нe嫆B��|}��;�>��I�gQ1%�p*"��Km���n�sC-��-�<M0��fe��ִ�%���
мE�Ӗ���v:d�$�&ᄾ`=�s�|����K)R�FI�o����:@+��r��xX%�r)�w�?���nĎb��v>��ݞ[��Y��No��IQ��v�e���r�XsgZ�m�s��v�8�]B��x"a��BaN/���� �!�����:��O�ˊ���a�HC�,\d��@�n[%�ʚ�bK�Z��\����f�8q ȃaXǜy�+R��`���-������p��׉�!�@�.`4����e�O�d>i�;�T4s �qe@Ng�b2����#�4� 3�;�7�~iz�@�)�.:$X+G0�-����`�%g�&�֐��(Ӥ��3խ��״^{Qժ�#��3��9�/�jBT��v���ƕL�|��.�-?b�:��V�t#N)�3�K?��f_[ nL�
{O1`C���j;K��:`���vB�N�?-�i�x_LM��؜
g�hs_`
USP��꽂��2.�G��t���o��@��_!��A,hM�	xG�@9�\�|��\�͚ݝB=QJ����K�NBF�C�f�4���@g.q�7�9��@�ȋp\Ow�A,|���1I�1@�{3���7!�d��:�����G�3B���K���������U�d����c ����G���
��מۚ��X�t�$���%�34(Dس�U[k����:u��/�? �R�m�.�RazGn�<K���]C��t�G��F_||��g`�H�/�i;�4&V���-D�R^�l�y�h#��І�;�0��x_a1�k�M���.r�`����S�v84����_ ڞ`�eNC���Rkc��O��c�������Y{�ZӔ3zʘ�,�QJ!��C�δn��2)q.�j�憭���	po��L@�8���W��yJ{ӱD0��]�$� A��� A{;���5�q�`��Fh�jN�Zcy'}(8Pmqz���k"Huͤ�m��������W6!��ρ�ȃ����K��l��)�dLm\�կ@"��Sd!���,�=.`���O��f>.��f�t�S��U�P�Y蠾0�Kyg���/�?�"���o��⭦��+ťϰ�qe�X{�Z}t�݊f.e�)Eғ�������~pu�iFIMo���		�(��&kE�2��
�١$naL��eu��q`��l�A�͇]u�F2C�U����7�6��1��咋�)g�2{�9v�D��tQ�q�o�x|O�9�mC邯uz���.)5g�Z��OO����9�3�4H*$�m�'/��sq�[/0�8�O	��~]�o{GdӍ�U����/:Q��e��A��$cg��&L�#�co������o�H3 s��L�#7�o:<ou:��������ꫦ���C����N$,����iW��� �����u��4j5�f�;I�UN_�,v�P|P��T�����p_��ZGҖ�����#��� ���e�Wp|׿� 'F����Ȝ*4�{�zr�mi�s]q%`���>]p�Vp��Xh<�X�R�u�E�}�0f8�>uCʐ*9�X�iN4u�`�q�E�o���!8H������R~u4n0@qH���\-�<�d#&b�B�E�8a�S�����fQ�	Ȣ ������3�/��r��G��)�-�c]n�r��zv�4#��Sj�O>p�R=�>��w��F�R]����>�Rv��x��%Y=��.]MLq/oP5������K��~�$���uZ��S9�0����_4h՚��M���:���[����yĿ����d�Ğe���N���$��@�:~��ͤ���Z����[|n�Ѱ1
`��߭�݈�q0}����ܽnpl����0���B�7d��p�'�ƩV���Y�xTc奫2�%�"���@0C��L���������<~�f��g���V[�?����\�@�-4�q}�z�1f1G2�p��S(��7�|R$��$p�P��Q;╃Q,!�`�C��2�A�_��>QxWK������}�8*i#�TPL��V$��{
	V ��
~}V�*?�X��܊?	�����ͯ�����C�7T�p���u�\�e������=���x�;
^� B���+2��s���k`���@X-d�8t�>Oo�,�%�j� �����0o��I�D��JM��A	[Ar��AF�a<�]@��g6�`4����8% ���޴)!����G��DVxS��E�d��%Bi�ҏخ�a558�G�	����ѳ
�YE�4��!���p�w;�݁N�S����-��J:a��ͅ_
�f#k�T W��}kmЩ�����V{���0t�e�c�����i�G͓�9�n�EŅ�	l�u�������`��?_ׅ���)s;oM�0��hJO�	�p��az�&}�N�u ��ō�y\xW��-������n��o
:�A� =ц"rx�1)]�|U�p�0pL��J��������M��±�8c��z=,�~��N5��5�#�qO�ljUM��ʘ;W �	}h��v�M��(����wwQMb�f�Q�!],üj]�S*�y����H@��M����,���D���Ne�س�p5A����O����P��]�K�����J�I�V�9i���k�	(��v�C�T�M@H��N�Ņ��rx���g�"�Ix  N����!UJ��L�2���6ZCi��$�,�������'���UCprۅh�e`���G3���bL�˱�F����X╹����}��2�q� A}�!�J[��d"���1��;���R���%X?���|b�зcM	1m%ڤʽ��7���Ιt���1o���=Hpzz�"�>� ��+ϋy�F!�æ�\�R�֌��x�<C�~��
�%$��	!�W�Aa���2��2�؛D�L4���Of���B���HBo/ȇ�@U5[=P��I<��8���y`�(
o�pwD'��2�/�;���z
�_)Y�i�W|ă����V�ƚ��m��lo�F	�09���uN~ee(5!j�I�zFAr]�G�ޯ�Yȫ�#�Qu�8U���"j���SF;��p`�t�Q�J��ҳ��T<\���(�6�A�X���:��I�Ĳ$��( (�h�� ��c;%8���%FT�*���xW|j�@��TWܗ��B��Et!���tC�,��dO������Z�xJ�ި_?e�書��N>֏4��u�~W�h����,v_�T�`I["i[�2v�W?=�K*0@],�Y���)��� �t��\���w1Xl�Z�Xr�T��JM���$М*�|�E"�g�7r�4�E��_��aڥ��t��o�<P������%��>ؙ.{�_"�L�����JJ z���C��{���*�BS>��x���7X�G�6H��`� P��C�}RQ�/�@������a��-�b$�i�D.�x�e8uW���SbE��zeį1o���䅞��u��G�+�>eR��ӶV>�t����<�[L�1���;�gm;n��hT�$�p`]�|�o�ݱ�yy ��i4� ,|.4cnX�����ͷ�a��b��­�Cm��ə���J�w�$�u��J�`�,/�⾛���El<��Ȼ�0�1�h�u����ӏ-6��M�qH��0q<�=��5����
��n���1�_]3�_��:1��CS|p��"�^�M�^�[��+ע��
g �n�H�lm-5�� )%|��CF�vx��1�3�'J+q8�3K�V=�PF�!Fz�rV�L �ֱ/"zk��cؕ]��W���ರڠ�_=�<Kt3��i�]���,��'e)X46��+�a��(0~X�EF��y4�i����v�/Iu�Hl�@��6��#��̪M��<3��kj!,��x3!V����J~���q��d�O+��F��j�/� �U~��tj�a��҃�&o?i�M�q@����kCt����s���Ё��G��t��N�&�5FM՞ϸd'�����Y�Z�]�N_� �AqR���
�N?({�����&�B+���C���L�p0����D�枇��61�%Zx��tR&��ֶun��U�l�'m����~���u������E�d�T�� �S'���3	'e���� �y����V�-|}C�/Ou�B�aQFb��
a���������\yȂх�kf�/�\�����;��9!ӓ [��`4�]c� ���A�ND|�"8�t7���u لQ�`"�Ϯ��w�!�@����h�T[H�:�=G`�rq��i��*G;�O�8~+�i�4��H���dWm��Ԑ�&}�^Z���̛L���=��a����:-��7㿊C6P�>=�4'T�t�z��@0��k���0`�,V,���r��F"%�?�uV4|R���;Z*���ަдn��lz,��-<�ߎp��z���ԅ��1���g�u/����C�"$�#K�x1#p� b~��m��W�9)Q/
���l=���r[��Y2��j>��?J�V���Y�0���ܒ�+.�����R"#�l�o���?�����eh��o���Dn��]E�
���t�Z�@�X�8���G��Z�Ң���+�0�w��~G������k����s��O9�+�5�&��k<���gA[%漮�g��^��p�E�r��?86Q�� ��EJc.��f.��-�CVc�D�a�߹��_����x^��_N�0,�N��(m|ߜ
�1e���JN�Z��hu����}& �*� ȣR�l�x��A&�$	HO�� �f��.uY���2H=���i��z���bV�+���g��7�cl�9�8L��S2P�A�O��=�
�.�Ch�Ń�9��$������^��H��埇�J߾Mh\t��^}q �ʛ�30%Xq$1���	�n���5i�3;�s����o�݁1��)���nw��D� ;�]�ؠ����ڼ��������P��1��5��u"ЂF��m�<Y"��p����4h&�T�J���k۩Ўv��6Bʲ	Sm����|NS'�=��.�v��}K.#0��)y�Ο*x��!��kU�&cf�^�W�\�9��7A���:t���%�c�"'�k�BXa8�R��]��>zR',?fˇ�ޝ7��ؓ-z7�0JV{�����ƅ�}����P��d�n��A��vn���ox�[COƂ&���y����[�;|���i��v����F������e22�t���.j���@"A8�hp�tG��,��7o���ѫ�D��^�AB��C����:�?vJ�%Q(%�@�ߢiR���	{����(������Cք�v�}�ɝ�Pǐ[q��'$���[�\��`��dP��jqp��5_�,ζ��E��i&���^n�4εx檁p��kUԁ�U�A��r!����"vq�F�E�>�PN�1�l:$z��KǽW�&T"Q+޴&���n�@�l�k�AAu�����Ǐuq1H6��S�%%<U�m�����O ��@��I0x�p�{��DW;9d�  0YL�A�D�+5��*�
�Oԟ����^nɟ�i�CA�A���)_e{�'t����j܂��pe�U���|� ��Ar�6=9A�2����,FL)�Ǿ�1�`�C�dЂ��δ�vY��Nq4̞A�p��-�HkW��:��\Oja'�
��	ѢTt��G�����vNR��G�49エp����lu�I�+���lC��	��.�b�،����zuQ>s�+/������Y���_��*s�r���>�+0�aȓ8AWL�ے 0�Q��5p�0�7�`�h2�y?"�3��#t#�v�D�E��3!��H��@���Z��2��q�n�Kqp$���~G��yz�\Z8E�f'p�uu�5A�
ԑ$��G��;bU`$z����VY�j9t�ȣk�#��v��I���Z�PT}`jvYS^1���P����#p��}N�GvC
�.��ﴙtti�ё�BL%��z/111����!�x����`3�Q�Ó���w�]*��E$x	o�i$,�֯ZH+Ou�r��b� ��s�=�⺅�/�Z�x�z.~I���@�[o�U�������8�L�og�}�ѭ��7%<��+��yV����^6C'F8�2<��Q�aP�&�����I�Y���t%����^�L%T���C_��zB�~�k��v���DV?����-w��I:.v���/�C��3�v�w�lx���{�k(m��1�Tf��S��}�>�4(�@Y�[T����3�<4ф�Ț��Yƕ���X��-m(b���p?H헗p�i�ֿ$��Z��O ezy�$��W�ck,S�5
�>ǥD�3�h�lYI��6k�%6�t�rY���0�I]L]��u$,���?XH�@s���Rl��8�Q6�w�R�{s Gjs�L����p���O~T�@��D��=R����/_Z6&�!;+f#&ٔ^�d��Dݱ�o�;t6?��	�CխȉT�R%ܩ�����:�?�j�3�T��ò�9Ya�MBb�~BY�^at�"�_Y�����Ô�*���fZ<4|�Q�9��#u���ʼ�'�?���<V.��י̈́�u
À�:�
r�Ag��	��7����A�6���(iŠA��ܧ�cb���;���Á���<�eG�{*ɘ8�K>���,�Kg�A����c%fʉe@���0
���*lӔ�8��ތ|O�ǉ˕u�cyab�F��O�@��$�h�D+�li�9���N�Ղ��� �q�g���c�8AJ��_�D�D�p-���Lm�CF'��Ѡ*�����3+m��`(��#�/A�T4��s�xMݐo��5����tKQ?s;rB�_�3��SQכs��� �4�tP�Z��4�*Q���<ѭp�K���PѠ��+"IJ��0F�/���O\�+���Pp�H��](lFߥ>6}Zɗ	v�تDu�U�(�������`�`;���\��X�O����_��F'M�?xFF���r���&�����:���As~ \�n��Mߪ��L���ţ��=��Z�s�d,k���n�,4G%�%o��}�!:{���UI#���ߜ �� �Ȝ����z��-a��6��D��8����G&�_2,�;���l�N��;9a`�g;N<G]�2�W n�����O0��(Xw�#�"U�����m���
�H�'��V�9�cE� >�F.�Ahc�(8#�PkW0��5���� .�\�mD�6�4���G�eI�:�Z���gzlY+��'��/ɑ�p},��*���
Pt�|�����\	��7���,X�b ���n��4�����V9�¥����go���B���� �Y�<v�'Ju�	!�*�f�֟�c�]�,�Y��U�����UT�iP"���=���
��4��SL�	�����Y���/}�ײ	ւA`�x�6d4���.�?�2�Ӈ�׿z����z~>���9��l���+���H������~��uQ��J�qȮ�1���#�܃�Бט L��s�rv�Csa�څMV?M����b�r�-�ŭ0�v�o<�w�~�J�}��JX�82��L饝��b��{�H.�����zP�UV7��ԎR�I$�99ٲ %4�_�wI������G�UN"� ����,�}��pi[iqH\��|�3I~ke�	��f�[XF	e�8D���W&N������ݿ?���:�q���	�p���~g�J]��Q�Y$��s�%��=n��r�B����{�W[��?��{��|�8����VF���e�I}>%�5���Ok�%�vc��7��׮ w]�M�!?j٢�f��ȸ�[`Z��A��(��˯㦴/Լ�͔8�-�>�ʢ�WK׎K>��db��LTvעG��jSW�S-�ࠋ���2Q��-��뵫�_���$C���`�1���x��gȩ�9���-�+<J��+��̓^��z��#х�3�	�>�ED�d\�#�1F�C2V�=Z��z�kw�`%jP�93Eru�a@�o>:}Z� ��a]o/����������ـR�6�&�A�Wğ(T�d�;��#x] �*'ih F��ȇf�Bc(�̕��o{1�U�R=Q�$�2	����HzCۺ��C��QR�	�/7�����q�A(�o�z�����)���u��l�JVTl��S�ۄ
�uʊ�O��mT[?� ���<�U�c�^���^s�*.`C�/Nن�y�Om+	�iI$�FՖG�dU��Gw\�����.�A�v��qk'��[�)B���A1�oZ�\�6���ˋ�����h��t����/c��=�7��K������0�y���g�ƙ�,�Ti� v����0p�Q���~�mI�����P|�#@����p'?kt�a�Ι��`aĊd?LՈ�7�]�(�T���w��Ɔ�����z��]�r�|e�������'	�������g�ʿ;�6�S���Û���ս> L���d�3�dr�)F�LZS=��Z�LƬy2��fE6�6%�25bD$+��b��!dp$�sB���y��yuD��j=�\:�
��|X@��<���aF���o��f�Y�I��}���>#]��� +����?�[��E���T�r��0��1���cYT�Z�M��v�=R%5�4}��f�y񙡁�����6@�7�|ӓ�h$rVUov=�H�2��Xo���F"�v�n�p�r~��*B �4�����|����`�x>{��� ���\�D}���#�K�:�;T����NCb}�tF}�@#+�,x�:Qa����G�u!.��3\꽹�_{S�5�F_�kχ���h5U�(]�o���a��x�����+3[IwAq�c��\�eL�m�5�spE����瓡�J�F�u%Y�p+�C�.F���LH���+����P����uu�1Ǻ3�1�1<�Z�	�6j�s�S5E�Y�#�����Ёa�}�S��A� ��'�_ޖ�Tu
��uw�����	�*7�i#��e�a}���l0�b��n��ؓ��RZ��$=zi+#��I ���.�<ՙ�[/�iO�M�n[И.M���;n���n|�9׶+�$�+s��3����C�*�������a�E����^���ڐ-�^����@����U���0�ܲ��'�1ʘ��@C�}N�L[��$�Ъ���H�B筑p�d����T�*6�.x��\QT���iݠ!4�O;�8��C�~�v 2�ÿ��P&���r����i���=f�������Y�7H&�Jj�ƍs�O�P��v��)��jaNT-!�L񎑘iOl�T[q��?	�(��U��6���ɰxL����"���j������%�1Q�Ӵ���9,I���4�IXe��̟���8 ��\pɏz�1 d���@��@$��-���Y�g f���v9Y��Li���0K�^��k"��j��"��\ɀ#�eVs�����[�g�ߞ�z��6H���
� �օ��ى;�{�Vu���]A�J����ڏ���r@x$���*]�d��9;ƛ������/N�]��O��&�@
*�pڦX�@&xJ�-A��aiLr�Y�fE>����QJ�9�7�z�!�+'X`�kQ��0�9�J�K��N������Iu�'rT �vi�@�؛D��"J��K�as�������J�Mj!�t�d��P �g�u��A�WI��M�l�/�ت�7�M���3�������n�P`w��Q1<�LD������ܺs������]l�k��P^���rg&7�R���6�w���]��4��`�
$i�6q�h 7�&	3N��ڴɍK|W����F,���B;T�H���g�'�����?.�O[�v/Ĵm[?�08=����srǜx��v����]m��Ƥy �+�1G����@��e
��	"O�Lm�MW:���U�,D�)��^sx�9�m��z���ng(M�J��Mo��~��)1������B���)��!���#�k@��Y:�?-C�h�� �W0% �0���O��<O�?k�W�d#D'�b8�!`�9�
3�}S0T|����|�5��9"���S}�G�\��jV
<��%�,��b�¶�p��j�b3��?�c�9�Gx� ��>E�u?KLq~_���/�V��hl�� ��Ai�X��[�Pq���Y��i_��`z��{���"��FMU�My�פ=����B���$�U`�dd��'1�_���m��A�j��;Nk��*?� ���������Z���Fy�鑲q!qw#H�7�<�+�c���7���AF:BCIb��!mt˯�K���չ!�׻�8���v�X�}�X|0����H b^n�|���Po�" QB�mwQ�ھ%i�|��>��V���	���l�O�z`�93��lY�EDT��K�;8-+�n%�'x�l=��y#R}�@���bG�(�]�2_�jI&�s�ì<��j�����C��>Al�b;��*�2��ߪثe�8ߵ^�G�9��]�4ѹ�gk���/� 1��F����b��R��t�im����b��F]�����].|t�/۠d�:L2��VJh.���K��jW0ԇ\�u@�͛~(O������8�� a���w�3����u������u2u|s: ;����P��?�Q�炊G8��.�1>8�(�Ꭹx�����A�PZ�	�C鴾�6WРw�Q۵�.�h���������ꊫ�ܿ-��͸Q^͋��_>�`�/�w&c��O���ù�ʾ�<TS��Оb�jsj�����%��7x�N*[
ɣ���"���7Έ���D����+�k�/�p�;�:� �ՎW�c܈#PPw��0���
V�4h�
�R~5H��8���2#Db�&�Mب@��&�fȋ}Z������\���>��dǣN��p���(�n��=<vT�V
�_�� ���6���ޅp鴼�Zc�_b�B�(���SG��K�<�>qi#'�4��$0iC��c��{= ��ؗ܇�iT��e�L��>!��c�h�_�����[1��o������\��,����;�;A����>�	^@��I�i7� ғq@'�m�8����p�{ :�=���Q@۪�'c�m�� �G�N���I~�<7$�wR�!�F����.���hYPm�9��������9D3�^������'��n�w78���:,�#B�~C����S��r�X������ˠ0Õ��/ܙ7g�݅�����?�22�<��TÚ���-�H��]��:�: ��Na�g[���ڽ���x���|(�A���;�����M�7K�X�ܛ;�;��B��h$�]�_`���%�=�=㹬���_���#�"j���c�ߗ��.��RO�!��*���&���o�+��v���ي��կhxu�������[�7�w ��o[�b"�C.����c5��H���6��4���NL��Z�`�"l��TN��mu֘t[�lF�*ֿ���ڥ�Cp �-�G�j.�;���[�5����Wu8Bs�G����`ϕ\k��E�U�3^�:�S��Z�9���Z>��(a�FG�e�mx�Q�YV;LW����+�n�HgY3�Xx�.�s$���#ATA�w)�D���U�H�ٻFQ����ѿ�� i�ߢ~"p3:���.
Q0��r$N��&����K���{J��AY[V�����eZ,�Ј1�}������3�^B$q5]�}T��j�й�n*�}-7��<��@ӕ�i����luC�$>�g�Ӄ��1u��vۀ�q ���e 
:$C�9�&�R��m�Q�m�l`F�+Ո�U�����tj<�i��GOKƼ���,'���,�r,#�2�����.�=�����+3M��l���%���xa`��w������o�1N�)�Ӑ�鳞]ߝ�~���./�9c?m�e|�ˈ��Ib~�ut>�~b@�l�Z"f*)y/�$lO��`p��P���Y���?;��X*��Yr�V�4 (�֞S�·���a�J�i����w���kc�Al��a09�=��fn�oSmO��~���@�ee^�����n����F�n��	�w}�Dح�@�&,�@h����ݲ6SV���	�}�����aY��ZH(('�ק�>-��~C�tx�Hūs�a�q�f �1��������[`���E�$~��#�3k�̡����=�3茯�aJ�P�d_���'r�2$
��O+U�D�L5�!i҅�T�s��h�v����;~�ȵa�,��\��Lk��2�K��-C6e4����`���j����1��S&�ٔ� hɁ��8p�W��1�~��OG_Ͳ�m��\�mu�DW�4�H�s�o�`1��������r�w]CT�C~t����b>߿���W�𜱈2�%����pbq�� ���km���{��y�$�߾{�'%�%2r�7Uᙦ���9�G{�g��=1�Ϊ��[�ĸ1v��?b�¹��J41�v	�x�����0T��1�U]��KC��"zS�2R8�Wg袖ƣ��߲q��پ)� �>#~|�c�)f���n����-�������χ�]�0����͍� ���-�u8�� �D��+�m j�dg�k���$���3H�o�p��&z���-j�����N�xO����pfS����l>
�鑆�t.ߩM���#WhQ����0���0w� �g��������8����9����
W�����ܵ/�m�yg��K ��'�F���/T�QZD$�壓hT�+��N0w*��r�g�[�����]�p��z@������/}�o���u��7����03�����}�ʟ�l}�7eW� 5`�'���J[B�o��f:k%��Ы����b�q��'�~�xkp���3��V�L8jnhO�K��CJ�=���-3�~�䁧��g(A4n�Jm�z�s�^��Cu��Ɩs_�N�9�|d�u,^Y�7%���`�G}:�eL~��f<���S�r��������2;<��4��	O	��:���3��WW��3񤾆�m�k��Y@�%\�h�+�a4r
��U�}��R�Z\��?��~���ݲ�3��7���j:>���k�JDkca�h���Ͷ�94�Dn-"}�o1��1��f�@�>d��" A>�ڑy㗔��x�J�53<�ܶ�K��D[(9��Bd`<�fȀz���yr���{F�������u̮R�� �m��+w5�+j�w��jdx{3����$��.��*�z5Z;�/�1�e����_�R�����A�w������}�uv�_��t=��V�
|�y����*�CaZ�e�K�UL������ޭ�!��Cn�l}�;�-MX$7�i��0���/W�j�8E`��{ށ��9�|㞙O��'�gE*�3�8���$�)g6&W�_�_�O�u"M1z�!Y�
��E��`,�D��4M�2�k3�c���^̀iwP�\�q�t"�����49w�P��)�Ʀ.�t̓k`���+C�懸�$�Mx�N@����A��β)��E_���N�2���b�Fj�21<Xy��`|�f��H������_�.�+?�ðr*�B���X�a��я�$cs�E��:�����a��ij�bn�јcU�uG|7宐/�+����U'�R; �i��Y����ʪ�XN���+��i��T������.�q*����׬�fm��}jռ��6 ��hu�XP��E�p;w��s���\`lVPW�m����)FH���A�|��G��7 !|��4ZZKP���&�) ~�fL1U9G�h���WE����(8(��� 4<�}H�������*c�ju[�^H�7�?e���L��J~,���}�{�H��8{��U!��zxGy~a��J��o����ф��Q9	)?/Z�;�}�@
�(H[�DZ̡�!���*����F�F�y>g)�
���-6pF�[Rq�C����jW)��O�U��%]'�T4Qeh���u�69����Aۻ��5����[��N~�4�ߘ@���P&�'��oӠ��40�����Aj`��Zv��@q�h���m=TM���M�_iD�sbu�6*��=ۇE�A�o�-��Nfg��Odz�t��Ot��Kb[<�$��0	=ddahBz�M��"�O�P[Q��x�L��"�;?+�ñ;�~n@+�������3j򛐱�xx��*���{u�l�Z ���J������v�:����W:�K��0R_��$�"� ��ӥ5�`������AS���3� ����A��=���:8(��E�۵����05ܶfH��U�����O���`,�o MF;	���zҁ	u����:0/�X�ȴp��W;5++�����c�l�.�����
.�(g�<�^`�B���!g���Vk���9�8�E2����	�<xx��If]w�w4����ÀWԂ��3�>�O ۸�	1S,�.���k�.)ɞu�F��k����(:��_��Z�SF[|��\XU����ZZ �陨��ַ�=�jl��~�MÆ2)G�-�W�\�
�Nt���D@ω�ZV}mlm�K�Л�k�&�ʧ@{3�N��sJFR���T�(]�<�j$DM��D&B#1�<�Y���K�]lJS��F@8�&ݤO8�-�,:`�
�z�y���o�B�������h��?���Z�{�ɞ*�!�
K�!����xD�SY��.}	��Q=������|U��jv�,���zt	I�.p�,�����0M�'^�{���O��Nÿ�P�����Y�K�&BQi�u/�P��Ѝ�0ŏ�Џ4t}L�1Tڑ5Lw�|�W���	�:�����S�����%\�^�Tᖉ���L8:2��4���Xk	����M0�ɤh���O�L�.$S�W�XZ��N	�i�،����L
J^� �������dT��O5+�E�´no;X�e�UE��_�W�7��t��1��q=������'�3�j��KB��f*��6Z��BgT�~��(� ���+���Z�Mq/;V������G$����u�G*�����F�Ӽ�G���(g�F�ʹPXš��ՙ����`��gn��g�L��&��EJ��}?ykv�}�+�Q�w�B�dc�<Eљ?�u��L4fY2y�j��c����̮L��X�,����k���	��F7԰
� �(�[��ŗ;ټu��}�M��1@���0ZcȜE[FN2�uP�����I<�b�G�:�Ըz��֘>����~�qY�W�z��ѿ�MXb�O��S
J d�A)�3�
��%����m�}�t�`$&S,n�nre�f��~��|:�Ƴz�w�ݓ|��z�L�?o�֓��!餜5��=��A29n��#"��p�$Bm^��ϳ���*Ӧ�TA�3s�6m�*��A��Τ,l���J�6�-�����[����ؑ�,�ҌW�Q�:_-vTf!�6	�U��V���\�_�a�V`d�;Gl)��['��6=*
�yS�'��T�����|9��o�[�+�E�i b�0�"/^t�'abt�^��X�0�]h F�W��������e�����w�P5�ϻ�we���,%����T�S.����ܜ���Ն�����G�/;�u�.�&��.����֒h��"���\{�˟n	%o�*D�?��An��,6��C�R�����W�\�Pg&�|NmZ�b������Qg)�m�i��>�f9�)o|��[ݙ��%Sb��l�n�f �����|����a~+2N���22�%S�qˈk�6$nΤ��m��
��@��뫒"ٯ�F@_b�u�
 7H��%�.�P��Dj����M�Q�k�����3x*Set�E)d���4w�#L���`E ��>X% I��ǥ��2��Ui�
=��kJ���E�w��0u����w�y��q0x[׶�mU������Ux��vwv���q���.�w����W��;n�@xr�1��E�"����@�ktZQ�����p�:�l��/���Y�â��'�U���\���٣+�(j~w�s�뺒�jq�X6�q)����BA�4���o�t��'�@���ۊ�Q��.�H�:���ڞ�;f���xQ��{�u���r�"N�ݟ{���B+�Bc|"��O����c��=f*&FU��Flx�QY^k�tu�-ٿ���)�ê��
w��t��"C/2�k���Ʒ݆f�V����R�g���u#G�7*�$��D���k_v��g��>_����U�ɞxF�yh��y��S���i�Ȥ��ov	/�~�r?b�,���^�!��Ln��5=ڍ՞��pp����N��
�5e֒��}r�B֝��Qi}ڮ�}/��~ߏ"�y�����Dkbl���N��3���i��wI������:ub�b�D�DH<a���M)���O����@��Fϒ3�	�TޱI`��/U3G�,�a�qtz�����v��z��e[&Ga�YQ�n獃]�{H�#j�P5�w2 #i����M��=��[}b���k�p���:"A����H���8�L?��||h�^��u3���a���B�Y���Sɰ4���'�TH���u��#N����F�˄����xv�����Ի��������˛����a�f1qE�9f�$�DU����(� ����%�&�s�"���&�|.�t��C�v@H�ipN�0IG]$ԵjaX3�n@�6d�R�k~H��c�]w�ݝ�#�
[��[K��b�Uс<�ę�p��@���z��d����1��
�H]&�R�w]���rn7���w>�W7K���8�1�� ��.�ו�N�䕓��&�S��{�F����.��5����n:�>_�����Ft��'�ek����B;�1��|�FA�W劂�wa�u�8�IHt<js�>�a�9�ɮ)����w}�
��7��탑�#�����%s-5_ո3��iHG�u�z�f��'ˢ��C�f=D���2l������.�=	��n����3>�DT���5XqɄ��9ki:�$��Z@ꢧ�t���{r�����
4�pO9�S��rF�rT�X�[�n�,IOX�Eg�qI^<�WвSb���Ϙ����So��<�ѣ���*���:�h�d�;��w�rջ��Ywce��6�9�����MOǛ�^ߦŻ�;�<(������/��Œg�C��Ƿ��,��H�C~��F��o�5i�梆=�=�ګ��e�c"3�4|�d�[����ѯ����y�{Je/�����$��t��7�v~9�yJ�Wgp�kF�z{�1�}�4]z�4�R�ظ�C�><9~�SF��
�8����b�0����� �R�)�1|�	��i�B'"�
/ ov��n��9H#ݏ����V����O��/���׃;u�	W��^�0=0A���A��6y��lv�`�������0���/{|�=9��t�h�V���;<�:c�8�jE1a�� �����z��+�-u�nw~��$�C��LϬ܊�����!��C�w"�3޽�����Q���h�Nx�͂p�XK��Q���8z�C?E���~{jZ���
�8��gC�W�b0��'�?H�?�uD���T�7�F�?m��o ����ϖ�9|F��f���1if'�&���Q���Z���ugn�rӗS-�i,��&8����Plaf_	����=���/�=5>�!��\I%��ȮnK2�x�eE1�b�M�xXuJ+� ��r��bb"��o�J?���碆�~[�t�����!���v��0�����%WB��c�(��S���'+��`w}�["U`-���{=���(&�sO�V9���xH3Cn�6m����")lf_3�c$#�u��
Ĵ�(�D�Kڽ1�e��u�^�|ki��1P�#�L%|�t��ezd�r���%iGtZ���II�k�v[��*d�f3��|i&��Sv��S_䆷�>�/e��5W���~tY�
�W�-��������0\�㡧�-�ʰ�g)3�!�%*�C{ú`�݈��ӻw�&*��7��Є��Q���Ѭi��?�z�MV]��CE�յX���S����`j��'П��z%i��,���L���<h���"���p�ǣb�k�t?�ّ��A;Z��RY2��=�$��ŉ�&����e'�ޒ6X���x�Ã�6��،=���܂�>^���V".Zx�\�/(���A�]�#����nYq����>��G��Kz+����y�^������67�֍	QM	*oʩ���Y�hu&�]�[���G����YJM��љ�n���`RNw������ݠE�?܁_�I<^:DG;��z�T�wg��Q�TGg:��\���;�#G7����i^�FͿ�Y
K|�p*�UBpv��iTQ��d^r����ûP����׼��{R{Ƿ�v�"���n�v_����_��ˑ9��@������ۮ��� I����>U���`.i������J(�Xd�]�&yE�I�n��e2c(��1;�.� h��7,�g���}���Z����r���Ec�x�}�qL$��`���	,�M�Z4Rm�����%&9/� ��21$3�xLf��/į-q@`�vK%�����Z�W�G�4�wJ/��G80ي�[%�`�co)8���ڛ%�_UN��@���Z{C�@���!UT�&2�_p��"�|�X�jzN i���{F�N[��*Q��-�7����3pu���3¤J5G����G�,c�wG@���g��Pߥ�,c�[y��l�FL
�A@C6�������$mI��Π�tL�,�B1�B6�
b���`/ó>,>!9Z�f�xz2!�~RWUF�<E �m1��/�G;�iW�j�8긓�$_\iU!�<o���@���&��nq �[�<�c�A4��⦐�|���3؈�	�)P�#x��i�rg�����=�'����c���8I�a��A-��/����f�d�	:K.L�a2�PT��s�޵��җ!:k�~$�J�%��Fj@�ƈ&���	����E�8r��o��^c�e��w|���z��6Sk��]��	J�iUD3�Y��� ;Q�{(~� 0F��]������k�qe�ev q�f=��Վ3n���)��u,@]&=jI[�X�4a;�٪�����7����}<��h��{��f����@V!��,)��9����fXf@Qb���d���L�n8�����m����?x.y�?�FKW��B�E��k3j.Y�Cw�m��S�N� �T����Kyqf��n���_+N̫�Xy��b�2Q�x�����x=Ϲ1,a���*��(gR!1��x؂_�BdeDְ�mbM��̵.1�,`���:1����D�ܕ�aH
���B�� ���Lh��%��0���睤oKi���k���Ns.E=�>8x���,${��/�KR�~Q{b8���cCM�[j1ِ�"w�c�#L���'2'$y?�#|4'�Ya���a�Ӟɏ7֍�zoe}1Ey��Ƃjz�����J+�ѐ� m���j3�W0Yb��S�I��ʐ�VYi/Z�CE,r��=<�E�~'��ڞ��7d�G��(��E^:p�pE��E�����B"��6m;��s�=M�<� w+�D|���p������_��1�)R��&P��(h&�8�|Cs�ƘJ�oh����>��L<<�e�Պ���$k�!ٟS�Q,E����,â�[�F2z�p:����SAiR�F���;��T�
Sx����2�jl�[c���$��bV�M&�$�o�iY��
����{(+&1�Z����O��Ӳ쏡
����.[BkT%�1��` �):)K��w9Q��Ɠ8_Q��ξ��a�GE�&Y`��s��WeG��<�aC����(���hiRsLi�$�ЛG���៥����< ��������{E�>��I�N��tX�ha����Z�͸�������\.X%�1��|����b��b}+���H�4��_r
V/<�Uv6�x��.T0
�z�C����r��A�^7ѷ�^�"��YA�3��޶�@�P��Wi�W	��^;em[�%�R���4�?a[���ocwf�xg���Q�+�U��.�M�Q,�F���n�$aB� �6�Y�?��^�iBW()����n����D�i\VTW^l7(��G2���Jx�d\�r�'Ѿ���^YJ�� 0�%�$>a^�ϛy]���P�=��8��=��7��)I(��L��oU!�M���s1� �@���+V���&2��$�)N1�G0��b|��Z��+�v}�B�������ETC������"�"^��F{�(�+4�o{Kk(=<<w�pR�(i|���%% ����82��sR�g|� 6%J������{���5�Tr�����(�(�B��-*�R���XK���]ٵ����jHj᷏�#t=�S]*F�4с�칊�tfư����� \]`�H�Z�]�o���W�A�i݁c,c]0��I���)EU���d��> �������*���|��?Xܛŋ���'�X�J�C�*��@)���s`fu�,�<�=�-�\k�&�%��Ӆ����� t��{۶![��oAx��NR�tr�J�;z�g�����@�P��t�}�A�JO�ٞm�0 ݍ�i�T(;��ܑK5��������*�d�*\Q$`�<D͹��f�M����='�k�S&���c�i�-JS�-g�˕{�Gg�#�f)܀����BnW�K��\�{��r��TIC�a_ș��m��^*�LJO�bo)2���T�x�/Ⱦn�!�i��� ���}��[���[��o��E�v��)��r�57�d�mⴳz�oE\J,�6��W��*���'�l��7�4d�$�����Y��r!��3���b�|3�_�;'d���k~@�g�t)��[� %����Wy&D�������`�yn2�4��>͏=�у����3 |�bכwο��?Ӯ�7��q��tfy�oe�sF�ث�b"[{���ٟȈ6�HQZ� �#��ܦ܀�ʿ|b��j��+���M�i]�i<�Yj�!��0�M��C��%3��rܗ � V&Q}j=`�f�`�}�qƻ��1rX0�&�i��O2؝�:�@�a���ֆr1�2���m��x伐�u��aHG^�g���}�ێO�E7ȏX�k��E��b��uY���_cpI|�xL
�e�]�w�o�z��[��L{q�ݎPRg�X<c���Ѝ�*��Ե^2�ϗo��,i�_��g1��w�<�,�xh�4��48��`��m�[����\�*�nH=��R��}9�_�ys(�'�g��+5�P��p���ؔr���l��c�Oo*�1�-���"�ĳ #�#��e�=��+i��|
h���%t\vfU��Xj6�ACy��Ba��!T�_˺�����Z�lǼ@�9�Q��@�`,�!�@�ɟDi̖/��?���oQ0�Z�"�z�o�̈ݛ�p��G��g�h��P���6�� ��s�'c�h�i�7���ф�(��?��5���frJ�
uO��S`6�pJ2��6;�ʰ�q �k�]UO;�X�#���=������`k���G	�o��P�"voHqސ��ۖ ���M7n�{����R�6D쌠$Z�5�j�#w񼈰����?�vU��	��K#M�%��5EU���`� ��~���S�ɚ�U�����gޣ��X��X��_O%�(3ϊ�5����]�TZ��ز�Q`��^�R�Ӱ�nEb���/��#�������I�V�w�^�c�O�~v���\��7�aSM�g�'��E.�ʶ�& ؘ������;.�8��Js[ȏ��3��=������Z�´��ɘ�z�߰ݤ.YU��N��<�M��_�r�J@�+�]���%���b�2�VC����t�S���Á�
�~n���H�������g7<r;F1�nٕ����Q��Y��$�����pG �� I��N�W9ߓ��O\�����Ta�{x�D��od	��F���i�q�cEߒ�R֎���1�����ˤU3������F��p��Y�����!��m�n�����J6�������z��F]�D:u!4�4B�ܶt˗x� ��������Hōx紬1�<pCby��S�J��3��Q(�,k�̚�%Q�$�oΡ�C��1��]V�nX��H��cRh1���c�W�옐/����}e^ ��}uO�^�}��IX�U;��Ȋ������c���~�Ǘ- �l8��u�`/�^\$��C*$1���E �sG�6'S�&J�I��ٖAJrV�
�R0�u`q,����A�%b�)[Bؑ�n`uC��˞��*�K�.�g�ޮ_%�$�bY�}� ~��PB��^HZ��A�B�]li6�z{%m_�{ַ�Ѡb\ė��c�~�����̟xP�8��H~�U�z�K�����X��ݛ��K��[���d�M�%��Z�s;���Y�'�Dr������+��� ��{����u��0�e�03TY��֥��։�a�����%@�#�^^�>��|x1ƪxP�Á+4��(�.��<���@K붌�#<�Ċx��oƯ.�[�1w�O�W9祻�l.�ȇב�OJ�^G���g`$�����V6:zCHʳD:�s�ҷvs�R#��&Sm�N׻��/L���'��Z�;�GlDx]/m�u�]�zlߟ{ύ+�.!0����%���gP��"��X-��3U�e�pwV1�Jxg1���ɠ���x��&6����g-����	/�-�~�Q�^
9�v~��=ۘ�g��|�� QR�b��X�?�ƃݸY˕W���t��P!������]��E���%R��_��>[��#��[�IO8��4#5И�9o�?��Zu�q0��.�v Z�>`�3/��ڸ	$t?�\wՂ~�bEpo�jQ�9Mq`����9w05ެi��1�0p\E7/�!�<>ܢPh��tw�6NY�@���0�^��Ϳ*d�i8#�y_�X��	�T?��t���_$�'r��A@�`�$��jy�n�vC����wu������W�3��=`��^�Ȣ&<������u�\�JX���[�?�;v�{�,���k��n��i	z�Q� 	��.Խt��%�����Կ˞���S*�"��RYS����5!r�� 1OJR�R�
�+���#��f3;4)���rϹ�h@��v�h���5k� ��?ܽ\���}��kNe��2����/�N�ԏ>��5Lj��ԧ��f�+V��f��כ���t�|�����c*ӕ��B&?���O!�ʎi%��F�2�;�,�C�R��B���#9�(��AySК���_x�b8����Wv�̩>��U�N�~�U�%[H��*K=9�F�GH�;�?���4(`�Fw�j��i�d����@�g����y���N}[cr��� 9�Aw��W������b3�w���h�;�u�>c~%��'A�$�+�4���[SMP�(��u�}*�{*�\��A��`{�?T���0փ�ZB�U3Y>3�f�9.pI~��fA��m��e����б������A��J}���J0�QT]Ae.��a5D%~Ͳ������z�\��*)eL~~fo%=;	���7��m
y*����-�=��9
�RX�ѲhfL	_�诬{z*��eLw�\'���\ }զܸø��~����6ʹA��Q�DM��Q�ډ{�!H����ᎰVu+�o��?�JFAm�s{�qn07�l7�������7܂PU{q���otXȦ��8�������H�;�i�ؘ����^��[v�W��aL�F2�d�����۶-=�zY��*��~^��ߧ��=��R7Fʀ��c����z�@,�ǩ�G�j����&o�1��+Оh�7�.A:Gވ�l����ѵ�)S}� ^�g:��S'Ok�:����h�H�~�'�u:��K %�o�bm��� ��t|����;�s:�s\�^;�ɻWf��.� ��ЊK#ò��#F �(��uL=75z
�g��0���ǒ��Y^�� )v�� �p£��N���Oh�A8	��_��,b�4L�����S� `� &R̎lv�gÕ����?�Ӡ����x���)���ъ���|�;�4�^	q'/�Dc��x�C!��r�ڃ �O��AJ)�غд�}�.�6O!vt��UL���CԀ���>���n�;��E,M�<����t��,hþ8d�,� ����ls�CI�dK�wu��f ���T��s���nY?7/w>�9�wp�ޗ��!I�,��
K�� �q5�׾OE��&�ř��3_Áp�hHY��N��D��k�'�o��~��Z���7�l�|���w�u,^
/�(��@ɝt<i�t௹�ob{gr-q�2������r��������2d�6]�]dԱ�ZK���_�����K��8mH�G�t�4���:!�bA�.Y>ǛE�ħWJ#c��U�������;�(b��ST�I���3��Ҁ�4����˺��_�̒7�V���+@h�bP��a�w: '���pk�w8�P���e/��#d/ h�����+��J�K8C؀�V����9넍�	ė�ʟ\��L����A�I]+�H��͜�n��J$F�y�R'�<*�o�9���0�\1~V�.d���g�ĝrCH��k�)���t����҄�窰�1"�<V�Ԉed�#��2ӹ@0lK�栗Ѹ���1��Z��3�;/^C|��_�?�o�G[t���\�/޸/�
wJ
u�$C��`r�[f@ɔ�)�d����A�TEP��pl,NV!��S�Q�E�Lɣ�����LR]��~!'�p:�>;it�餌X=*���wq]�s딧U��8�O܁	j�ϻɞ�QP.�T!��y�ȡr�,!��� ��}����4����m�RHu��B*�>�7u�7	�ES,���(�]2F8T�N��Wl]��a�׻�f&$����?»�:'����C�gj���3�t����}qw�.�����?��nȽ�[�8�f[�'�h�*#�`�U6j=��#�*���F}�ـinT�-8�V����3e#�QF6F��?6mĭ	 �X��f	�wKj���^z���8�V��Y���3���V�d�'+z�:���u�;�Y�i�ą�����ʎ���.g���p6(�e�a�n�Y\8������X�T
�rDp�j��-hN �E|2���f�|jX&A�u�7�V���!�Ańa�8K/��4(`�5����0ڜg��u8�����?�ސX�|�u�hr ( ����{���9�qK�_gza��uCSA�2��V�W�Yr��>P�rY������~��۴��	h�ki�Ca+?y��T�� Y8�D|	���ot�<ً;d� |3��I��(�^��s�T��p[ǥ8�X�[���Օ���������H%B�z;;�bꛣd9Qy�*�j�1�ef�Q{=×��M��&�l
G�習H�*�64ԛ�T�o���ɸTLj@�XZBR־��J��#��u;b�K9T��m\i�h0NF�Z�Xll�wo�w|>Qғ�?^�Bi��!B����V��,���eA�1w���*Z�B�<ǒ��{���Ω�؇C��i��W3�5�%X�V��$���mX�&_�-w>�&t��g�ZM!�9#���x!�l���j�F1!}��扳���#���Bʬs{��Ik��Ud� KmB�כ��-Z�t6�p�������F�@@Q-�&�%T�+މ���Q��U-sz���0GR����q���*��ώ#���t}�'��(w2�	WAs
)Nny�"�$�C�6*7(ᮧ�MŲ[���<�C�ORb(�ʵ&��[S�_:�Ӥ�*H���U�-س���p�U�	�5��p*p*9�(�� N��G��P=���&�z��w�T�ep|YP
�P�v=� (�8q��Hw+`�����x�lo����K�	��Z��J�}��ol� ��g��0�)glV�����aM��hG����S�DZ^��bA�/���9c��>�}g��d�W����1�buC=D6�^E��r� fTH1��u5@�G[��Ɔ���ۊ��It�lѮ:_��5��k�8~.�>&l��z����[�S �<{��u?�3����| ��0�a���ކ�Y?�xG?* �Z�%,��̷�������3&�c���~��Ӑ�Q?~����y��qxAֆ2X�D�fn�����n�>
�I�J���r�EtY�g��KQ9�롎����&Y�C��(�PH��&�!8\=�T�k&d�X�s�R-�pM�ş��S��,�ZŨd���O�%ه��c�E��61�rN�r ����dDڵ�������J�l�,�f�o?l�
|� b�^��14�58w��-Y�����x����8�`��r�Y�9>	5�9r��.Z���Ʌ�o�Q���J2D�vG+ߠPTMF���S�H�^��g�0�8�ےL����ˌ���!�)9�����U>U��?��&���.v���Sm%�����v�$���Yv�������T�u�g���D��������
A���v%yE���KX�fE��٪�G���Y�Q��@D��$3�O��n�)��w�Ew�H@q�T��5+1/9����i&<�y��C@@sv�6C�}d����I�v@�k�	���5Xզ�T�Ă�Q=�a���1���4��L �ŭ%P���$�M��jx��$����>ͤ������`�i��^�O�0��7�`������p+�(^�[>F�ko�t�Ac�K�V�Vl�8T�Ewgb��2:9��F	�8YP����*Z��^,�(��LZ&Bv�S>DC��"˔�*9�@�К���n�j6}��hh�l5N�@ˊ�URL�s�wr�`��X�t���T����:V3��x�}@e�Մ�h��kX�G ���[�of��R��y��I�.adY �6Tڳ3R�(�
8�) ���g'Ϯ�&��;�ܸ��w�r�W���1���ȧ�b���}�����P����O����|:����	HĠʿ���"~W��OJ��F�+�9�L����!�+X ���-e~������å&�*OӜ΍�©א7�I�x�36�-�Zn$�{py�V�s���q7��Lu�z�ȵ�|���T�Ew���]��&U�p�w��{-�����y��ܸ1i�����9Z��1���$��{�ׇ�TFa������7�)]w���=��QA�,�_z����^�"��<s��ٙ;QP�c��s�oN���q���a]a.s/�1MW�d�'��gc��_���_�B�і1��؟����'Y�,������mn.�sLL&޷�
���qJЏYg�CqW%�x����֖�цn%��%gPd�O�^?��]N;�W/����7�P��y㕬�����z u}-!���x�z�:�Ϸ������%`�(����背����(��7(����`q�٠e!��9�q'�����;��s"IRfX��ނ��D5��5cJ�	H�Cpm$ʪ���F� ;y����Y�1R��]ʻq�X�K� _��x�M�}v�<7����Ph��gG�=ol�yR�!4&�t8��`�(>R���6��>oAC�>4k|���
� #Jx-� ������Æʈ����J��&=�v"#ΤY���ҥ�Ui��͉J�������\x��Ȳ��F|��yR�f��?�B�)�e�����ކ+��hY85�ߚs�cB��w�V¼R�7\1i��	�����>Y���Q70<����ku&:[�/�B��s��|������'��a�Gё�a��N�ᤄ�h�z�a<�@.bs;��Į jd�η�c맆�'�����'Ȩ�5�9��؏�F}�?�H�,}1���V�d(��������=>A5��:)�;� ƀfi�k��:X^���S���ܪP���y��"�]�\쐢�}όF����2�U0��� �޶����t��Nر�1�+�N�NVx��2; �٪\�4��'�ǚ�'�bh�*M������Ya$��gwCw��X��L�b#W	
�{�8Re(��*����z
�����&Pj��D=�:�����W���z%��(TK�^ђu��[��c{(D�9�s���w�$�@�^9�̜��-"֤!�K3@i_箚���בi�"�)�(9 қ���>A��Tc�oY�����7'Ж��
��L��"���0p�I�*�\�O�`G�]�8����q�7�n��E���@4��O�!ƙ��h��;�� ���f�2f�(��i�+�d�x�-���p��yz�=����܂nQ"�G��r��9�^3)jM�_���++�_|z�B��$�=��FiZ�F�I�� �tZh�+u�{4c�A�n*��}����~�3����i�_i)��BR�Vzx.�>R.w��7�P<���1�}uȌ�;Dn�=����w���ZFu�U.�W1���@@�(<2�ڙ9��!�p`>F�_y�Y?z��E�~U��:�L��I�S����	�	���s���f�:s3/p�����QR���()X�U#������M���}�2;"r�P��(=)9�.~�;@6Wh��/qZ���'v��9�v�s����[WkK��$"���!S��A	:�N�H-�=(��B"�{���Ͼ���(��	�Q�4��h��̼�jm ���CwlW������D$,~��oX�,��O��?��3�jʧ������A�k����q����$��X�E��x��Ϋ�>i���f��\��5���oO��'a���n38:4K=`����8�>۽���JE�2�(g<��fp���s�Hp@�OGS{����z#�u�X�t�<��B�{��84 �i`���BW�G�j��נ��`�b��h1�1�����|#��.B:��lZ7P�,��sY�Ni��(��ՁL�,�F=�P���o@�����}�%��`)���b:j��5��6��������Cjr*�%�
�?p�֏Ì�)b�H*}����j�:)�Մ��C{]��������3amp��Vq��_��#�(>г�9�P�h�(���ZvI������|��`���BR��������H';��S���p�:?���=U����*e�Q��uo뭜X���"��c�kE"�1��~���{6���W5�`��ex��?�k9n�e�8 tW��ky2���}Yl�[h)�����B����N�����ߓ���ͩB<V�E{1X��b���d`�UἪ2���'_w]b���k�Ʉz�7�<3���Ir�ʔSDUv"v㦕�1�a=}��gEl�{4y���C�7�Noψ%���s�V=��e���pֶW���-~�3gx�5u*.�ձ��í� �
�J��RCHt���#�(i�~Ϛ�Q�F6K�����_7Q��f�A���3s�����}��Z��Z��/�-���M6�E��V׿�y��|�-���͏���)�J�/����d͸!x�P��%��d��4�;�^�D
Y�r��t�J	��I^?t�t-�L}i5x�ܬ]|�KS�v6i*7�0��\B��w���}�8 �q=p!�Pԑ��U�Z�U�����r��~�r��А�@$N0�qC����H�V���'k,&пE��/eJf
�%1���P��t���w@=(n����g�<S3��h�v;�Y�Qئ�����m���(#����A@/��c�"���ͮ��k��Չݦ� �pX��o�1��ب�C	�x�9)�P1@��?���G��I�n��N��;z�&�+����:�fS��U/ �/d�'��E �:9k����O��M�N"h"L���ϴ��Z6����&U���`hT�e�=������U����/�f���K�4�� t�x8Lp9�?uJ�z�̬�3�7�pB�ʸ������ί�(�2�X+���P�O�=&��c�����hby?�p�M�ݡ^[�,]���	��ƪ�6�N>�S��s4V�� �޲v25�Z���n�%�[/�F�qi��#,<!��˟������`
�蝻Ff�8�Y��`��X�VΪ���\4"��B�;����_��Q��ʨܝؾ�� p:���Ƕ�_��_ZQ�2��B�m��ACF.�Y��
`l����$�+J���H!A��$�k��p���u�A����@��q���V�p$1�b:�/JfY?���k��&��` ��t缜�������U�gp�>A�T�������\��g��+��.�V;�X�Aa/�=��p3�8E~g�גc���v ��:Q�&��]A�����07��m���Q'&n	B�^3�Ӏk�XB��-p}A$LzE�ժE��ފ�@�hi�
�> ~z���_^�Hl>��pa��R���b�{�f*�k<O>�׭k8�h�u�����F�䶿�k`����5�ߺ1�6�f���:-9<>;���'���7;��q�M:�*�TM���T!�.6�=%^yܓI���u.x��ҋsZ3e��"e����"�jn+��R���8�c�[%�k:��ԏ�i�4�(Kє9�UAɁP̉��
ш�ޟ��rI��?{Wc�GI���;@OSΪ
�=y��rt"��A1z���	����"��N�,"�J��-��U�KMy0�w ���#�7�}�����cx�!��Mω�!a�{� ���X:f�.������ !�� �.I�x�:�.�~�Uη[)k�2���TƱ�n:c��ٟ��! �煑��X2��8՜��1��,'�R|R0��OS�4�7�O�Cq���6|A��lS�������%An� u;rC$�W�"�}a<7-���8)��e��Y���֪:ti�1�M'��1�_~�PC�~_�
H������QrZ��Oݴ
{/� wR�D�3]�l��q����e�P;̥nZ%�wc
���L��_�ü�%��;)HZ��ƥ]C
Oۆ�x��)# �<����>t&Z_Lw��h�%k]=�O�'���,���3N����r�l��zkU�<����6�!L8�t׊d��'�]73Co�^n'���N����8f�t��簥+�Z����5������p�=w�2x�.�]�lJ�V ����
D��q�#�A+]� �e.�=��|禮AQ����m#��2��,�wN����`M��x��o����T�$��t��@�|j����k˩��!W�0H_7�/E6�����I�2	�if�-\��>�0t�EX���ŷG���b�����Y@oY���JMc'27�Pk�џ�W�)�� ���3�w�@yNtv�q��N ��U��"��l���,�.��c��L1Μ5GD�^X;q��9�EƷ���T^M��_�KDgv�pQH+"�V�`璀w��U���b�;i�Ft�p�����k/pM����� E��ϐ�ɳ� ��d�܃��eb%u N���v�~K}1��Ι�ЇyAr'U�R��sjog�A�~��GW
��e߾�@U�͎��bg�o�����SXғR����E%vr��2��U&�FC��+�u=����ob=6�ʒ'������R������X��8	��j��x	�w!���Y[z�ɤ{|ګΛ^��T5=YT���k�?��{op	Yi��"���}:s�!�=aOɚi���g9`y��3l��XC ��G<�,�!;�api?�Hխ������v�?J�Pt_��sO� t>m�r:�n�K)$��.7M��nZ��Ze��/[e_���:��C��U� ^���E�$'������"�� ��Ӯ����2/>?��7)�S�oD
�{}��{`ZԎ?�h�ˑ��P�ȷ�I�"�Q%�G*Mܾ��8�R( ZL�!��0���ZgEB���KJ�߫ϸ�p�z�R�	�ڊ��/����SНu�F�s��Wo�H�{A�)$sN����+����S�����Ѡp�R�bCf�z�"����XK��'#��*i�!%2�Z9%�u�������:��|^�2b��L��a�+J��f[���c������z􄰬�F�86��:q�����p�TiIpM���q��b鉠��,�-�� 
�������2�#�C�� O�����҇L����r�춟��'x	���q�KG��.��|z�M@�ôzuπ��ļ���Foe5V�3b�Q�l*�c	��~�A�����r2a�<�R}�o>W��"l���0�f�	��N�!$+��r��W!�n&�E�#<���%� ���f�N�M��U����Y��Y�t�#�T�6��-:t}S��&����03�Dʸ���i�e[��L'���nي�c*[���ó6���.����q���r��{^�+>=CM/��c�͞��go܂lۏ	�f�xl}_���]2ME���n��b�MLV���I��xN^.6����=�Kf�������ל�|O~<jͷVo�r?���4+��T0+�5�*��
����n�dH�`}j=���tF
π~��Rg� :�Hh�޺���Ŏ�Fl��U��P���W^�s��e�M�!/���G�v럯����~�Z�8Lf�v�%�m���,c��Z�M<�w}z�i>w�e動v�������$:vf��Su۟����[:1�L�����	��eځu��_����;ΰ�m���u���hS�� "j�t��~~_9�ob�r��o'Z���������2K_J�n�Ξb�HA�~AӼ��zzϺ��Y[�{'�]���i�.��2e瘥�
��:�2��oJ�F\��a$6BƱ�.1-��+`B�c&���5�eU��>��%o��K(Y��{�+n?�N��`������s�l���s�|��n����n�5clr���P/Q���ӕ�l����/.�Q�N=q7�},���eU ������{ʹ�"�~�10�����F
mye��.�@�z��s���x�o��g�v[V��Q!�Gu���Z��om�V��AҮs׏��w���3�H����UR߃ީcl���H� 1�"e��L�Z�Q&e�5Cu�06yj�Z��W\��?��?���r^-�ݮa��I-��1�#�ns�ƈ�ӳ�P9���(0)�=���F+.eR�P�M��ӣ�˷{�&�Bu֊�o�R�H���Ru��h�+�Ss�Q �����Z��7j��誘0կ�č��jI�	��i���1��~Z�� �J�ގ�_��4ʒ�=68!5h=s���w`��I� �:DE���1{l_	<�7L�pYF��,h��'@�i%���oB���~VU9qf2ά�Tm��f&oF�.�}���v�����/b��ZF؄�;vW9g��Y�i]�lo����ޖ�0G�&�ѽ�qD���O����r�
\H��V���y=HMz�]����]^��D��d�" "�����6��&U�
�e���{Wg�3����G�5(i�G/��!��mw5��_Il���y�`�δX�v�3w93Z�S/t�a�Nɜ{L�X_�s��OE&�B��;��8g�g���)�prY�+�3�ŭ��q�}�7�]J�g���S��@�E܎��V�~��M�r;��Ti���>�����Lz���C��,�
�C��uɘ����M#�_�`�!�$ ڒ3�5����Đc��#�Q?����H ����E�2�,����.&d��{���[��a&8E;�REJ���8*�l�'K�Q�����+�}X�l	l�j4���� �\�?�O�~�<u�<�@%/i�����l�m�tZ�Jm���&þ�]�@׷���Y5�3��5��k!�����_�DB,�l��$aA�[�l�꾎t��U7�!`J��/����AS]Q�L�7�a5���7<��N�Ӿ�����W`�J���W3A��
�	�!�ƌ�X�q�ܪ����=�+ע������TZ�P%}]h�ߺ��ȸ��:��xg�>�����*��lyE˟=���tUeF��/�M]�>�rt�D��.Q�8����_r��S�B̠qf�[�CU��쥧9B'�_�ܠ>0=��xZ@P@��吕�6�V[LėjnMs���q8����noj���e��t�T/�I��Q���ڵk���J.@�VH�3�n57��j)o�*B��Z�
���D�ĩS���t����KJ�D�h0��u��8�����9Y�!���Zm>��=P\~�'W����Id,���ْ���H�"tl�*yԎd�m��������L>&]�K��0Hm�C�FC��k��ʫ6���jrƬ1�
�C8��R������`���AФX*�i��g��5.�`kG�7P�|>CC��m�ڌu/���8�l��8�r��� ��c����v����y�UR�lO����Ȧm/W���B��|��������|or�PP�G���l!i�N3�̱<��*�L�]eC�\��7#Q��EX�ʱ��׏�b�����O5��i+�UV��`(���=��&	���B�Q_;c���kʤ>��/
k��(�Р��>�� ��ֿ/WT�73�&�N �@:�mx Ζ'=%�^�?|3rx�|XA�����)���1����(k:�-��#e~O��=�+�1��3�\���Q�3
�!�V��DA������i���ly#.Ѿ�/�tт�Z'�s�J����ϔF�"����������ٜ��Ș�<V#���Qe����W�2/���w54y~��=���v�5mdSh��K��7إ�<�qԶt�ѐJ�N��k�p-�k8D��L�iI��D����n5�X#���H` ���߫pS�ѽ�f�����&�~A:��G'F毎����gO���%����ݩ���^�"��l�� NX���z���D��c���GzN�vod�|�Tv������r�q���)��a�����A3zR.��̴�����`�����r�[0:&	�w(�����sp<c��-n��Ȟ�x����**��"cd<y��@�g�.�\B;� E���DYd���5Sii�DUy[�_�<��4�˃�'}/թR'D��r�i3�����!HAG��~��e�I���!�#/Q�3!�P�2�����Z���|c��Lp��*�:v4�A��58Q�l�����}�}u�����2]�����P0�W���ز=e{�� !|����
��
4�hY+��y��b����^�q<��_4��q��S�`����_h���+�c ��z�2S���������S��g�����m��T�aX�M�ڛT�g~�	�x�n���� eQ�nh��XJ?֫��fc�2����1J����[����
�0Ȃ-t��փ���0�����M,DZ�\ѿ�����:�
m����+z�!��>�ź�����*r=��S3c�.X5�yw�_ -��_���2�U�i|/y[{i�_��N2��cS�OԻ�����#��f���f0���B�x5�L��i�2D44
^((�f�Oÿq4e�W[�6&Q�A�8b�	eD��x��@~�29��k��eo�K$������JN��@��b�ჁL��GZj�ZdD�K=?�M��8rJ;`�Ilńu�����i|�ǐ��e��B���/MN0_L���$27�΃
�

VK��w:�h�c#\r�:��Ǹ������o�J��	�% ��H_���7���ɡmWP��F��J{�a+Cv�� G��Rs�ٜ��W��#O����!��H���0��ʱ�I��;�s$��B�o�B�!иƢq��A�˸%�/g�-����[F5���|�虴���XL��<S�,�~H޹����p'꾬 ��_�\�ny�����4��lD5ِ8�WaU��K�%yG#����|L 4�A�lL�̖��Lܷ�)N���։v!X�!@�܉,��5��W��h��M����FP��.CG>�o(@	f��c!%��ҿ@����+*H�q����{&�@��1��Q����2���.��dE�ʽ�ލ��[����Om��ዾ�r�N�\�(!E���g�:I�O%�B5�~���8�m���K5�M�+�k�ۦѩ{'@�_J�pDD�+��H�c���u����n��'��(e�m~��)���@�����u�̓6r5|�h���٬�H�W/���C���qoeH�I�KM��+��KuH�ƍ��� f�����i�<��*���\��>V*�ى��I�e�~މ
�@�m�X�<N2F��o�U�G�
|k�ۃ��	9��C@̑���qb9��y�
N��7��Ѻ���AD!���(U�,/Q�C�k��R�yٌ�3Fс�1E_�]��Z%���k���}Cn�+�V�w��vx�W}sJ�q�z�'�l�@4�
�mz4�|�z-v8z��mД������}U�k��_�6CQ��Y����+�=���HAzx���O	'��Ք�$Yo���-r���±%l)]a��0C�Wqr�K�l]M��R�EF������K%sɌt�{�#���_\�0���{;�:�W�.����"k��}�vذ��1�����Vˉ�&@���1�����7z02��B�#����5`�M��W�6(鶼>�����~�K.��-J�K�^���Oi,D���؛�����Ĥ����Q��t�@�
�o��@������Ȩ2�o>�c�U"��a1��vؼ�#�"n��v�K�
�G�9�Km󧁇��W0�~	4?�%ps�$��)G�(��	�)��E�u�TȂߔ'bnJ�zP���+O�Ԣy?�o>W�G�Τ��l����ʽ�S�gL���^���J`6��<��u03�"�;��nԄa��.R0�~���N�؁//��M.6�S;f7��r/��y$jCrv`�n����˞�.1�[H3F˕F.���I��bp�a^�ޔsl�Xl�9���L�!׆HT@���������!`G4�^���-���	�#W/W��1ܥH�~��d�/�����G����$�x��p��v_v4����sJ���:�-zz$����� �ǉ[�L��ڤt������( �
͑_M2�V�X^�UD�{"����*�W��6��.������W^�*�b��c���P؏T�9l[������_�K�ObL�*�rpQ�L�+i}�Eώ|�>COW����F\��i9�~ �+0O@�c]��=lL�9��Eox�Lk��I�*��F�5cwZy��f��ߐG���Ԡ�K���}��n��ɡHo�}�{ԮN�.�u�|�������)�Z��L�'��/�@���-f�R�d�L,<�lP��ӱ�KXY5�S-= �NS�6Fg /~{�9���R�.��X��+N�؜Y�/����Rrؼo��e��&��-L|�(z��+�H	�\;��a���˽���z)�\��~֝Y�#�wF�{���u�lp�A��	�����!3��e�̑�JdȔj�vӘ�lۏm���~ ��i�_S�brT�����<P��$��{���!��gHI�[۪��BpW�=X�ECQ�d*��X��?�Hhx�|S׫ǋ�k*|�}aK!3YԒ�+ſ_]�溼�}$n���I�dְ�W|��F�>⬆f��&|��I�D4\F�Grl>����<w��>n˯qE��9 G��	:���{���1� �K��Q��L�pkb��E%y�6�dZE�-��(e�I�ݻh���Z�*��=V%�KN/�>DiV�h�o$�_�\ � J,��mx�N�\�H|0§�q��w6���u��D�9��3�KZ���\�R`�������\'Fo��U��p��*V��%"�/�����&� ާ�N����&�dF��5Ȧ�s�l?&�fP�a~�%�����2Y�c��1e�3u�k��0��s�<F�m�6�KyJ�J���������Vj��ɗ�*��\0�" i�n'�]�-�K*V�+�q����u-��2a!�$p��vp�a�i�6���A^�c��x�-��}��b��o0�I�pM�3Ã-j�y���TU?�+781�-k0�(͈�~0���s���,���~��y�?V��{7�C'&'�|��$_γ2Ҝi�0K�A`�y�����\��_�m|Kn���<EL<EQL���2�d�t:V���V'
36����s�������3]E��Ďٜ��ςfO�|g�=�P*��>�e�,���J
hU�����`M�MK;k��_�E�A؛Q}��̈́`���i$�]����5�^�����o5���=� ���=�3�Elg4�?#�ŷe�l�V뮖
�|ƥ^/�:},����g�m|Qː.q���k��rʉ���cwz�t�~��������#�mn��Fu�~�	�b+�#�B�=(g]}W8�S��t_��N���B��u����Q�ؒ~�T_�b��V��Ը��}۝�j�Dj^2�N"�b�,���P�{f����=� ��?�4�@sX�2������<����z�& ��3)܎�҉�>S-�*�˸�gc�^�D.��25Q�"��@�$�h� #��U�e�<���TN�` ���}�h�`��Cbut�_�.�,�I.+wi,�T�W��<�l�@�?tC�*����N��Z�"v�6�Iԇ�w`I�ĪZǜ����"�`Ӣ���������������S�^3�:�;L`2*o@��ŔX�΃�\�z�&B�s�m�n�Y�!PM��
G�&�/BH� DQ_�j39e�co��\��k����> �o��[B_�^iɵv�*��^��)� ���m�%d���!��Y��/���w���c�ĽW�X|2�>yz�\��(�IҲkr,mJ.4��$���r?b]��R,�?#�^����j���8�[���k�>�Ϩ���<���[u���?r�fj��<~�n��qݩ���z�)�<\���t'7��i��J��I �|0�I��6��Q,r��U�OXF1����Yw��w�D�Z�v�Mw �A���Q	U-�]���.��*%D͛��鼥��sa�
&C��Mٹ{�^��٤X�4 �*�w�UY6��+#����.L �ټ�5��{�>F���?���zo1J�sa�M�ڔ/An���\"�x�?�'��W�ΰr�Ç,!!��D�+�d�	f�H�� 6��2�=�����;"� dFF�t�:3j{�Yn�?����|�O1qQ`^�M�7?t�֙%���� �Nͬ�����,Psޢ��_��y�E�#r����Z�vaV��)�{j�G�e^Ikv��@֗�#6���j��0Uz�A�@'hh��2eۼ�����iH��D���=!3�ݯ2a���3�rnŲT�E�L[�m�^�~�6�I)f� �6-z����;��5W�r��c�����G���J�u6�˶|ȺTe߰`����y���j�U|�H
�����B�ȕ_�^=�>=*�@D��̖�s�8�}�r���4ȗE��j��X ��Yix9��r�B6[>H�ܨ����$������d黅2'��i&i;��F�i��;��-����s�k�{�yw�;���j��/�*/��A�i^&��y����- ԁ�`�j#4���P��	��ƌ{V�
���		h�9B�)ͣ^+�,�g���v$��E�s��Е����ꎛsa��x��#� �z�p�,݈n�o;��ԁJ�dx:� ��=�w"���_�cps��K�k��iۖ�g��d�Yd�=��p�ªg� ,SD��)����z���)�&^�M-ҕSHk�*�.+�U����)�Zb1�:��O�݃�f'dE�H��������l�&��JQ����f��-2��E�ܢ~��AТ�E��#���A�壩�e��%X��%!4o�	U���<���+L���>/��.�\���Tq�%���/��܎�=����F�n=����W�R5%��c���2/t�47�.�R���V{��B��&�'�{n��ǆ�{�/Rb�n���n0W�0D5"�}6���/��p��N	Rbx&�p}o�؟�_XٜKy,�K��'.J�]0<���1y�J�˫pP��L�Fű� �J'�����Y���e@��l�}
2k�!'�w�}tw�l�92�Y��� 嵭����i��}}7�4�yt� 41�ͭ�/�8C�*��+�k4�f�t"G���"�� �? �cF������7>"�-,dp9r��F�-k���J9�\}�P�+^��&���=��,-Q^S�t���[�
��w�d��y��Y��#Fѽ�����#?���^�	'?u��0NEVݵ�Ƽ�I�����@��q�z@���x�y��6�[��5VG�Q8d��AG!]�jؤ>2��l�Ed�5�ݱ�[CH�Ĵ{p a1�1$��Ė�%�ߜ�噀��-�����c�,����
�V��,��J�{J�3�3�@IP�f�9������K:����qyl'���AE�����3�~����'T�p#נz|��8�A"�O*ǈ���o���У[W�1���Z�+1�j�]t^ W�kl�I>�B-��%ޘ(.�$߭sN�~��];���>��t����t)��;e}NH�ӳw�v�1���1�ø�F��㱾�*q������� ��v������}��~��A�8s����~Y A�Jy�E&@8Fn��l2)�8]û��3��eP������M����^�_We���V��<��L�����l�"(�h2��=� ���*�s<n��3T���<�E4�c����>����.�/[�9!lD�/Ft&�~�f#lk�۲<-���U���e�:9�hK���������3�0�-�eW��e��XC l��t?�T��(}��SA��b9Q��6]o�����J�Q�0 95!�F1�BJ%w������RR8m� �r)tH�a1aS�9s�D� ����*P&�}���\9�������7��;��n3#H�9��k�͖��A�����~tVw��uqspJ��	��&�){���,� �y� ��ZY3n��9Q�g�m���A���
��E�FF��q�J������c��M+��f����&��M��Y���)�T����B/�C�d4����ɉ~ ����Oc���	�"gB&k��E�S^X�8�Uz4�Ȑ_̖`���T@+=�c/��N���I�M��5T5Y�Ϝn �%�smX����N��Ӆ���lJ���,;	{Aܱ��|n5��]Հv�C�{~����������0îm����.�d�B�7y	{r�B~~�(=.��
�
�O|:�-RWC_�cQ���И���<T(A�S$c��v�f?B$j_"�t`�^Y1~�����-=���!|>3����d��~�Uc��c�s�9���U��0}&���^[3�v��m\o]���0�.K����ئ6@ޙ)7��_[���`9I^� �7�׊�9��{��SGS���� �<���~���*��i�U��3ڰ��5�/o�{�9[\ �/��U��g6�R3�U��AހVG�:0AD]�%������oaf�-FU�*���]�y{��n�W�|o�׉�a�u������~a��G�݄�T�p�w���2���j�&����U����L��G3�+�[
���n?��E��ͅ��'�a7S䤞[�������Ү!�]���Y�E��A��g�?!��DY�ӰJ��� 1�vy2�&�w��S��i��KR:�Dٜ0WEB߄��L-T	���j֒Cܚ�Yp��7)[Ӱ�`��n12!���R���LX�i+<'Ҳph��_ٰ�y��V��R����<���{;T!�\x�%6#Z�mŒ�а���Ů��9q2���ҋ�~N!�u�R��4��A�Yq0��kJ�OޓҋP|��Yǲ�bo;n�d�+�a��A5>�Q�HXeZ-�*�m�h1�|O?|��N4d:�r�$�3$Zk����JF�̥�#�}y�:�*b�xr�W��p��k*-b�Dl�x���_Q�Ĥ��T�H9����_�5�~TЀ��<,'v�8e[���u��x�.�@�uP<��� *��Y�����\��P�&��9f����A���-r�VDX�N#[�A������%��� +�$h�s薖�E�v��[IJ
+�F��8T�-x��Y�/��9���%���4��(�<`q� �)G)��(��1���6؈ݦ�LD3�1�#�M�q;NO�^��.�A�Nb�Ib��--v�mH�s���a��g�s���@[�[�5�+�_�|d��l���A��</�c��%4&��+��Ar	�R.�Y�����,,)� ���A�Jv����F�����AY�u��!O����	J=���)7��d��y���ʤBZ�<�t!�d��h��ЄAN��VV�jo8F#��X�!�ϊ��8Ӧ��|M_������?2 �����D!G?����X�;��(�ɥQX�8�+�+�r�A$_��7�8�]�_�I���r���cq=v���N(���O���z�>KU+A�tgi\qzq-�bs�|K�+&M6�e (��~�zl���#e�@*x�U���%b��k��n�Y+��铞lq����W�-�=\��BĨ��֩L��ש��_a�R�p�;�f{�f�Ŀ��f����}�|g��$sF��퀽��g7˺�4�2��֨�9y�tgd���G�]�l�D/���["�~�2&����7���;�H1hA �PԼE8˵��	{�B���=ȓ[`��v���&1;2���Ȍoύ�Ҕ�4�S"�8��p(�Q��B���k<]*�+6r�J$��7���t�xg(
:��4RF��T�Pj���sO�Y�yԵFxz�������NX����.����z���|��hl��Tn��a��W�����f��������C�fH����F��IO�8O̚-�-`��r�	�5�&�� ��R�T�p��v�&/�1[?ǔ�X���q�����#dkQj`31)�cc;��J9~�][;���N[�;=Q!���56QP�PAVg*���7Y-4yo`g7
~�D[�|���RQ�y��B5�	y$-��saUt��^7<|�9]���iA�.��P:'�����tU�I��Ɏ��o�+��|�w�j����g8\�f�KX����z�o?V�ۘ�:��L�~.�L@�mIھ�>0t*�kа�uw\���?�x01�"ݫ	��#R$h�f�n�X�q����ފ}��]�_�Ë�b�__*����ƽf'�N��_����݌��{��"�+
:,��S`�@6�Șz��]�����y2���۷�T򱰸r�O��1�� f��Gj��6�V���iJ��Q��|&�'�������z+���n���;W4]�0���$R�o�M[�^���O�[!MR�l��ޗY���A�JPr!�M�SO[�1F<}`�ܫ��AMr����y�.{rw�NBYG?S�{Ƙ��d+�WH>L�O�c�s�'8����]x�L��)Wғ��7W�L0{�I�ޕ.��aN��W!5��F@�?�¯RZu�'���P9{��G�P{���֊J�-Z�2�c�C��b͖2K�<�3����@EXb0���|">A_�c\���Y�l�f[�K�a�������2�4za��4���lh|S�4����ASy�seW��TY<�/i�%�a�	�@���d�f�\��@>z5p�?���"V;<��Xg�I ���O����ꇌ՗�a���AD�;yT;��nf���m�d�~����8�	����!!R�©a���6�`�a�;�`����t�n����_K��R災�e��� c��k�&Ot�k�峦�x�<na,4�D�ׂ<j1ᵃms�|���|ҷ��X�͊�.D�cJ��<WB:��_Q�qj��M}�^��u9]�5�w�Cr��2�Ś�ǭ�Խ���<Pa�Yn�+���g�*��L!�s�A��2 ������٧ͥq?�՝���q�~�	cˊ�7��C|�]���B��ɥ-�*�w���~��>mIӾ�i�M�4Wӝ�)�K�g�D���됆Rn�um������( &���m@o �!�;ZY����a�%��\���6��i��>�42H`N������ɞ��L ���\�;�(A㸁n���`N�+19(�,�<Y���6�B,.8��m <�i��^J���Bz�>������o��,0��k�W-�/p���}w�zǻ��@l������A�H�ԇ����V�D�Hl{�NA�o ;rWA��!}c�|�K�x�	xS5�1�ϲ"c)z�7Y��J8]_�m�L�Q����A*��>wI�� u��-�5|��.E��K4����T��5�8��^K-� �;�����ċT&*�J=�֍�<ys7��t�c��N(\
�?d{���S�¤2^x�'v%)�ag��⣡�<���Մm�Rb�l8�K�g7���"Y��Sy������8IƗ��1I��� ��=��Wu��=Ѥ����b懽(�A83�����:{��]��Z�ɖ���V��5�Ąn��F��������#�#��r�I��;���˴�W��Ƀ�Q�@�;�H1+��z:0j�R�(cy��+�6~�?(����
$��l�(�+ڀ&`���3/G�P�i�� �<���� H@)�?�CX�Җ���xK��HD:\
��M��A���F	����&2��4֮Cr�<D
�K.�hB��'������5�9�au5Qf�V���!���Ê����3���R�:rмcv���������? ͖I�T�%F�fowI5/�@�.�=����72_�Q
��|�\t��d�0�� �io/,>l������@
���晵�:�To�����3��"�c��6*,��q��x�Y���xypf��i���`O����Q�*/�Eެ�_� (2Z�P<)G�Ұ��5V�#0;�����(��C�����!��SH��1*oΡbbϹHULY��F��I���#4�trϾ.wm}_���].�	\��F����To)��x��"�0ꛋxtk�[�c���ouX8�C��XV�e�V흇��S(7p�-���<��������Qr���RM���젾�M���!z6̈́~X�����f�͇5�v�{����� ����-�U�7Q_\n��H�7;<�°�,cJ�ƅ�_����l��`NZH���l����P�Z&5��_i�m��R���gP'� uA�Β̚K迆�WD��J�l�b!���L��öq��^�_	稜�D[=ΝӅ}�l��P�hkww�9�1]g�e�'[��z/!����ď<e6�}��/�QS.�5�@.��,??3#�S|q�v�f���
F���\��q���b�$�I���34�pV����0��sS&�	0@0 S4~�3~F�I`�ʡ�:��k��ˏy��[�����ga&#^�RS��W�s��A�7D$sj��-#=��m
gf{�� Ǥ���$}s1x�oN/��L��3PlD̄MGf��@1:T�P���d{��*T����EK�ZSę3R�h�� ^_�L~����_}��0�q1Y�n��i@jF�)�fQ4$���N~��R�h`��7:�to1^U���S���M�G�<E�����^Ӑ�LQ�(=�9�T����+TŃI�_�l�m�F+��aE�3n*��&����ci�)Mp �O��m�PK��y��\[!k}ZfZ�<M�� ���gn&l��Z�ƞ'��u� �K�`,���f��k�������x����(�xQ.�˨���?����r�t�� �3���R��JR��B��b��D�
"$f�N��.����g ���ŝ�]J��"��K����H:�Ey �#�	O�J�F~P�P���=[��B�^�?��hЯ����)��C� px0$W	�<g�n��yaC$���11ve��+���01t�[����j� �Kv�.�(�j=]���E�'���q��T�=��){�08�j���Y{Jo���L��I�nڱ��G�Af^�a�v�DM}몑9S�}�ӡ�(�.붤f�n,z?ܟ4�6�%�?��(Al�g�\��s}O�ȆWUe��It3Bϰ�,h�k�����Y/JM��»;K��-c-2}��KKt�C��,�|�? p$v��MR;��d��7ݖГ߳fnw���b������c�@�05uemOx�V����dIgz�Vd�A��?�}K�;+�I̐H���r�x�M���b�ix��5�r,�z���;��\r�,�SV] CA���2�x�#Rn�<d�j��qm�G�-UՁ�	�ʤ7u�t��	:�Nn��+�t5�ᔤҮ�%�h5d�@m� لH����t�S�2�D��c��Y���X��W������z1�y��ƥ̮��n�?٬��t�ԟXE����� �U�x�:@���2�|�xR��Ҫ����p�����+�l�TU���~^�k�䅴�qs���	d�ۤ�&�ئ�y�~��$}�M�e}L�V���}V°�����*�$T�m������'��VO�g��|���|�?z^�" _r؟'٭usS���e�LE�!����f�2���l��V��Yp|���,�Ip�ֺ�XwO$F�a���`�����%m��s�ޭ��C�N��x����f�$^�|N5�NT�������D弈�.��!-����P`��s�	�''��h� �]����Ԧ��\r����K��/����t&�cN}B�zBM���"�|\&��~cN���4�Ռ��=3Ʈd���-��~DD$��Q�7��"��(y�\4���n�L�v*֚��ϵB�@m9;�^l���`�-S=���;.P ��!t������5��N�h,
������t�(]c2�����WŪ8Z�0�W���db�A
O����~X�O��Z*PY~����	�ۜ��r�@`$�n\exy�SWEw�խ&[]t%���Z��2��/ԕ����V�q�����q�צ,.׸��!1���j�;��_[�=`�ʹ�?J:<���yg3��j='^��m����0~&����jnl4�8s�?�Q����E�L�k�W�d�-�`@*�*:�b&�ˍ0&n0�D����xƺj*��RG�?�����) ��$tF^<��|��h���3e��NX#oW����B,�Fș�Cl�ݦ\�x[��p	��E'O�V�}���X�|_�b�?j�}��/h�{A�~�NR'w��@�B�����=�g��ك��'�֔H��F %�$ͭr�˚� �n����wd�HB��0-L�Zr�g��)�$�ٙ�b�?byP�*Cu����WA�� ʦ�P"��\ƪ�mD�vWd(�����\d_�:.g[+.���'.>�����ON\naT�$���~B����k�#�nB&\���i�/,��� �O�Y�enO��ז ����	c�{O~��ܯ�&�j����,��V6/����m'wQ�Ә�EV���M���d���OK���q谄��R�24Pz[R��m���D���sU��v���������Ԭ!\��y�{��ʔ��Q�πh��0���6?�Y�mK�L��d"����l|�mG�fH����n}"��*��r�@����q�����DY�&�d+�D�H�Ʒ�wL6G�Iz$��A߻�,7��&��u�uxHt��m������5�鵾�4�Y�zJ��U��ı/\���n�O��`�A
��IR�	�-�V]3��Ը^��\�����n��������:y�i���B�X�j���V߷3�&]9�r8:)�B��U��^ 39�	ٔ�<��QC�U���KxH���y�e��-LXv2Ǚ�S� ��R?-��S'��(D�MB�A�Tu���g���J?��jĘ���q�7	�a�����A�ʂ5����c�$pF�4Jx��9��R�tB�{OE6��0�Ð��E�-ڞ�Q�#� �W��u1����+I �q����\��@YR�Uj�I�!]k\��� 2��
�/�?��c�|ZM�TBB�ߣ���?����j�@�A��q�8�&�Y�ђ�s��{l}����{�KLuG1���Z���&��Lb<����/�P��m�{�� �*Pz���}�\�{m��=�.jU���w�����$ ��:	tw�m�������K��*+e�Y����G��buuK���b��n�Ӽ�O��V{:i`�ˡ�D�8Ltǣ�nX�N.C�i�SێMI��d����� ��v%�rdvYtF�ܵ���v���?$s�)l�Xo�W�`��T�}��7�f��-+uR<�.iK�s�\���z�~�s͵��Gd�#���A��jtWn�gS���)uH]?F�/Ӽ���9�=����p��99�����*s;(O�V�AZ>��J���5�1f#ELl�hӺ�����i��Һ��� ��DR,�.�ʔx�{�F=ٮ�`�A�=�I���O�r�����/eƕ��aټ[����r�Ӥ-B�|��:�*Z�p���V;�'��Yl`dC��t�؞��;���,A�k���&G<�Ȍ�"�2dD�8�F<�b�8u��� 7s���я��+ɲ��:���Ka7V@�{���'��!�}���p�b�~:/MF*w8����V,��+�s����Bv�ko�d�0l����h႔�)���?'�x䃡 � Q�'~�J=1U�.�y?���\�1��z)ӓN���,��h�aB|�Ǜ$Ci���ڡ�l���BN�p�����&���BDþP�F�^�ȧ%f�.p��#�p�'lfu���3Ez���6۵Ek�E�#z�i��ů�_f���ϣ�%��ޅv�C"0��'�x<� ��Z�=k���'G2�s��b|�S�V��߈N>vHl��=E1J�(!Ț��Ƕd��%ǰ$�&[▸�Y��|�R<����߬��7>��쬘n�xjH�%`�h��%3E�i��ѩ��{���=����"@I�����ohX�^F��7><[�4�&�>0G-y��N��&�̱?�z8���)�>˵׿.���!�W_T�K��	8ၻ�br���.��s��vb�����y��1RB2�� ?��˄5C�E5��T�UyY��M;�Hi̤����bY�e�ڗ0"��7㍺T.������'� ���xY�8&�H�C��xs��P�V*PZ��]�J��Z*�β�� ���V���4�1B_m��@�%MܬK�5�3����&��	��1�d],��CK���/��٭7�~+�q������L;US��܂���x�b���u�^h�6;GmA���@Z��
�2�DlU�r��8n���ygh���fL7汋��ZnP�g������$��b��+���{V[gXv�u�a���s�1m6K�iO�7���^� Ӳ޲����#L���d��xcN��$�^u�;�,�';��,�+��.G�x�� ��G���m�}����Ő�ا|��e������mkIQ�郷3ur��@�YcR󽔹�4�O�_��̀�k>�C�{���u�����¾��_�鄘��X��|K�*�z�<<�&E��3�"�.2�(}k���錴��+�ـaT�:͸W,.��[�l޺����	pd	8m�k �f�:��{���dbLj3�x����(�m~�J�xU��G���A�4I�@�M��kv���ˊ�Ё?�����Lɏ��ҷѫ?/��*y�y5�<n��(js��i�0�ϊAJ��#Y��b��
������
+�7hj�3��f��i3
�b#	M^�P,�)�$����Qt���@� �T���:��!B�����Ȋcu��{���	H�#]K~Ϲ��b��}�/�ճY���M�b9��[�(��Ϣ�����F��%���*�Շ=!R��r�m�_�!�-�_��6�+X
Ӈ��7�;D����JJa-]�����W�F"�?mF�U�mu�g�����|��Ce�)��^�;�±%�xmqz���~��ꑳL_���HV�x�if�9���>��p赣�##���s��2�k���0����F��O"׻ذ�+�H��ݻ��z�*0�n��|�x�Y�/k�����E�S%n�@�$�'#]W9�w��9��s�v���K�%��..�&�ȿ��v�^������џ�ȋ���W�NM#�xq��]��h&�(cP��hI�>tX���)Չŵ-W���B�⒔�.E���tfS�N�_(�1H	�q�����pK=��ހfx+������/���(T�@�q�� �F��b)�j�hs�Z�q[��	�-�Ӏ�w�B@�r2m�~��phl^�ޅ}�LD	���c٘	�o�[���&5Y�<&w�\0@�����!Q4�y{|3�p�H\�ܲ��Y_�;ߍ�1�5��؇�a�SQag"ߔ�,r���G3�<����?�?�!Z�?�M��2<v�Ӄ��9 �~���Q�B��<e�W�^�
,2/��c�˽�rP�=H�p�`8�ʁp�����h,��s�&���gݴ��l��d�����)��C$�'~n�n1��P	G_��a���Hvs)
 ���Q{�����V�� o�C�R�f\*H�U�����|��䄦_�,����Җ���5��=�B|���>����7��r8`/'6���R��2��׈>=-}a�
)o�f6V�P�b(K�vx��Uw�J���ɣ�B�j�E�����s��[u>�g�d<�0[�s4�B��Dӭ�#M��q��Q��(%�`E�����[ݓ�R���{��9#��DK���2��dͭ��q�(�'�:'��֨�t�[T��r%�"��X�?�k4\o��>k���+�@�Y�O�y:��IKKj��g�����I+�NG�����q����Ml"�m���y+L�KL��˭��Ȼ;�R�c�xK�n�"؈y--�7R�g3�O+ 	i�׃�
H�����-�1��W�h��:p�ɭK|�WghVz^͑dq���rf�2������q��"
�3kl&�/��n��Zz�I�cb�q���xf�F b'@�]�Mܛ�J��^0ȅGO��p4���&��H5�\9v/��C]�	K��x�RSa:�� �`|�E��By�T	:���m�=t���{��;����u�TPf>-�{�I�W+��x�G��`��E�e<y�S�(�id�AR9��?^#Lu��̏!H!Uv׮rL��Δ'�:[�pK�I���U�Yv��/�Xo&� ���>�Һ�,A�^�JiA*�Fn���+�H84�46��P-Q����j�Wy�E"�$�o�q�~��W���f��)��|�(X�����@���� ��;����W�� �A@Ā��#NP��-���8�=��1��ˏ2yё=g�{F��&D�j�Y�d��Ώ:k�3��T�V'��As�S�ߧ�IB�L����P5��Z}�+�QU�PL�ǈ8�Pu�-�Q�~)���\�d��5���b�'m��ȓ4e `Ńd����l�6����*1��^�,�m���	F���\2013ĹIڹQj�p�e���==�+�iu��c�1��2�Ǧ�õ�ckh��ݯÞ]�L^h���(yo��� �1]o#�5��e��U�qmF��Ȥ`�n}��c�3~�̇�zJ���W���Yo���1óPk��zȣ��P��~�z�O�������[�
��]��6�^�|x �ND���2	P���_G�Wؘq����wfU;��'9�*qf��`���V�
u������u�2������������ӊ��w��Kg�H�9H��l�H�d�0FXA�J0m��q����Ç$]b��������yB�.xa���o�@�\qH�뛲�{���p��:&�_q*Ey�J�Ȁ�RA�,��S˟��^��\[��q��T�\�\6�� eM�p>(���  �����$�-N;Hǜ�jk�w\\��ӽ�nP_7��EEq���/�|�r~,�?ov���æ�O�6t�f0&;Ǿ���KkQlc�/y 7�BW^�ǩs�gl�$����g(����ZF\b4��X�J�JE�������D� �beN]@�f,��9����4 ω���>UV��;��P%��h$O��3��a���<��w�r�+���hZ���l�t��q��%VĊ�?LAC� �y:�7�^ނ�����E=R��,�����&�2����6��F��iSg��, 1ޤH���u�
��ݖE�,M���F�%�n�����Ճ��11�������L��QҀE�aJ�����������pR��TB
K��b	�Ew�3��Z�J�"���.��Y�B�Ggӱ�$)���%u�Ǵ�|v����!I��b%M��K���A�*�/�hkݩ���g��;�����U��/u�F��E��D�v^-�?�b2b��J@��I��Ip�bͨHC���E��رi��0�����y�j���fOW#d�\�+*�P�on�3�y|a��M�O�2��[�t�a	f�/]���'�D)�/ׁ"p�>r��B�K
u@���q�{��k���Ah���'����*���'ا�$��;nSю�����,W!_�X��� ��f��җw�WZ?�T�ɋ%r�T(����*�C���)37�VP;�t��A�(���Y����h���B����A��ݿX�o:�A�.\<dn�_�E�����6��K����^�xj�YϸC~�|u%%�K��P�K�桨�1D]��1�'4O(��V]OU{7��9�9s�(�p==&L����3y�����A�����1�9�xKgn�����_'�)���FPD�9�NB
WZ�/R�����̫to�L|�5��:3!uc߼M��2��w�6�8�Յ�c��l�S��p��S�Om��{�\�S[��5�4U�j�sG�����wAg��8M�G�T�ϑ̫!�m�Yz���x\�نApl|4��R�=�+B�<��R�Ũ�AJ���qB�8|$ʜ���X�ID���}�G�I��ow<�Y�?�0��Y�%	0=��%�i�=�9.�5_�=�U�������R���'pSE�y~��ڿ��Bl��(9�g 
��Ѥ��:ˁ�M����3�&F�K��5�+�B��5s�bU'�="�ս������vN}.ﶛ�"!��#�r�f�q?�=2񑻏�/}]uv.R%�':V���Z���;��4�.�ԋ,��`��:���-ڗ$f:���y�Gőcܤ���P^�F�</mE��z�����y2OK��{"1w�/�U��m���Ǹ$�	�~��@���kѺ�����M��rR�� k��*)-�������|�7՜hԶcv�E ZT��ˏa��ƴ�r�w��ꢉKD/�4��u��~mk���|A�p��hH$�j����j�	C2�푶�Z��i����s6�*�g�V�CѷE���c�T�ܾɓ�\��MY��fq{�3���[Ⱥ�Q3\���)��o��
MӁ�`�ۤ��L�>�����	(��~l�6�^V��)��x���Ź�����d*�����CsN�j;2n=�+p�5$��s�C0�BZaإ����-�q���ȳ��W�WA"����ݘF��Ԍ�I)�E�2��H�~���Aj8����r���8P������ǚ���sŋv�ʱ�9C��oF
����#Ė��i��`7?F�'�[y�	�e�W�Ӥ"Ҏ;�(�Vyn6�f9�T��P��;?��������o�_c�Ŋ��IE�F%2%��0š�WYs.2vYM�ژ�=�$,4"΋eZ��#P<(-�%���#�w��{��ii�6֋P�}����U|��R�E�4!�Q��[(��a*c�2v���E&�]��N0��[s��r��ݑ���h��>G�[�|P�Q��Q��1�kM��]W	��K��Q)gF#�����5��|�V��w��*���-X��N��+' ؀"D��i�$�8��a���������+��Lc���g��5"�i����o���M���qn�n�Q�(T��G�C�R4ԓ�wSOBu�<;��q1=��{�@��c "��D*�s���M�/�����uBⴶ�~� ���.@�xVb�V���!HpLA�DH���d�� %L;����8����/���3|G
��c���?Mn?bZ]��t?q�ظx����;�B�-�c����Yk�I�ĩ��k��6�����;_Y�o���l}ꂼ�b���J͹���t�{v�r��u�����qG� �=�����:�@�T3�����yT�,��<S+�s7S�VFr�4�k�-A�|ۉ���!Mkm��u�&�@TJ���+�뗽���L����]�H�DQ��������P�gsB@N��eN���g�z�\�l���!�sm�I��i�˰=B!Ki	�
Y�:C-�nN�̝�c��H�&"�B ��QG	���z�O��
��B&�U4�/�ªM(�rM�2G�C�]��H^��;�΍~׫JX�̫(�����3���	���0�j	H h>ĵ&�����]2�t@A��{.?O���g�)s���#A���}��^ly4���Oq�)i�+����v�4�䐉���-j��o�Ȣ��I��D2	�gI.]C^�tⴓqs�*s\n��+0�W���n.�V
�B��_�q�8ɏ���=���OS��Ӱ}@'v͵`�+]�+�p��9�U��SM��q����K����|t���)Q2��Y9�ݵ�e�|�m�1mR`r'�/c�nî�|�[�.�8�kV���!L�r�u �����|`��^��~p�\����|�L��*b������YN�a��R��`
ֲLʢ�1��P�o<�K9��C��ӎ�U����^q�h.§}�-;OU��ȚT�Z�cR��-�	5�h��8VI&�9le�����R~�˙^�Ֆ������^@�0���8	ȫ;���-FN|e�f�@�c��x+	?�kG�Hh�H�5rE�̃5z��;~\QdTΦ��>�	Ð⟈� �#3^���a
�`f��l'��R�SN���29>�7�8h�v&��N�K�]��.��޿�cѾQN�1�*�Xȇq��K������@K�tRo�~s�>�N��%��������{��]�ڴ͠ō���V0Td]n
6M�)�U��	Y���z��v�Fg9���k��̘�
M���|�ÿ��01�M����:��۸��!���?�~���_W!�E��9_Y�ȸ߬�{PE���� �T9����ӫ}67�WT���3�7�vo׫A:ZOO;�w���ˇ���{jki��f�`S�������0�ϸ�M��㭭�"�/?B5V�������0i�M4f۱	H�* )�j��;M%�?,��>�ڛ���Vgr���7���v<�zX	�@d�����C��5e�g\�}n�^��<�Җ�4�����Iɦ-�R�!0N#�0�d���͝�������
3�bְ��'��w�ѵ".ۘ�j�1y��k�9�}U��bŕz'O��{�-��]㈀�j-��{�PT�m+�i1S�HB����ų��LC��,�&.Qi��M��C]k����g8�
rO�2���c��>�bd��i<a4o�|	�,��*Ka�BaտU�>�?8�I�a�O��}S]�kbZ����W�3��<5� &��N���oO���1�˙r�zu�>{�#�������u��u��5">�S�Y��.C!byf�u$!��k�.�<�����eY��ŷ<���O��8֪�ѱܶ���	�x��Ԝ#�& sΑ�"D#>g�r:G�$R@��h9\D�����- T����SV���Z�72��#>���|�BX�Ȁ�		���Os��d�:1YTD��L���I���f���@"�S��)��$ģ9W�T��j&�
bM!�}��W\�k�B~���	�|�\�v`@'���~	����$��6p�,L�~���F��!a�.{��@�_�N��}47|Lj��B�����;�]�ã7i�=n�tFw��ķ���@)F��5��^�������lPFp�5�N�+N�l>T�=f��P�+�%�XS�����}Y�@�A�?��c����`���欸�?GwOM�(H�<�)����V6���Ǧ��)Ĳ�X7�(RՂ)��z��S���98|�7����^�

���$��t��vr�M�Y�*��yNx?YJ��F�X@��Іg0��:�AHh�p�ǣDdL9o�={{�i��� �D����k���Wog���*�I��V�o��U�q�G
V���N��͍Ɉ�?�Iwu�W	з��y��
�� *\r�>���c^sO��-�����au����j�r
�i�S���^F�ṱ�C"����.:9Һyy_���0h��
v3�F'��̔�?g�VQ����aE��.�����ŐnF.&������!���"N�"9����f�/�Y(#7�Є̢���(�9�p���"d_w��,�Q�dog�2L��?(�RѬRK��]y�����h���%
�O���:�\�3D�h�_�tZڲ��Y��Q���e�Nȯ�\P-d���Z4|���}c�ߣ)<�sc7�=F�S�����8�~ 믓P�i��}����4��Sê��T�q9������}̿��W3�N�j�(�۾����vvCc;�=���'��j;�<j̏;��"U�u�r�Շ�6�b���fm�
@�-�+��X9�(tn�r0�nY]����Z3�����Q�t����`�V�� �(�T�|��v�o]��2k�ad�ڻx��FX�d�+Ÿ�MKр���aB�C�k�fzH9^��@��RCE�=�"�q�&�OO�}94{���i9a����]�"=د���
�=�6�bDX�;�c�ߞ� _�> B��vҐ�j�������|��� �[�k���w���t���)�h;�hx�6�>�o���6��^Cв �H�7ڇ�
�hb�^@��/:��r�	��@r�`���� ���w?ͺ`��7��Z������7�V��֭G�Z� |^d�@b���߶7������VC峻ڳ�@`�3Z�P�딪��]_b��4�_���*n��U��%�m#@q���Ha�������Z�rai�eB�9�w���5�%,�LIH�ql\u\�*%Cwеh;>6@��`���ڊYпZ��*㾦���B:إj%��	JO炪
14L<_��!�0�"�G�D0�<��^J��Ms��eo�iY^d���m�{�#�^��h.��]";�.EW����X���h+�D��^������o���c-��g�(��#)�g���=?������%� _�R�>Ql$�ME~;�C�l�&�Iz}^�	x���$V.c#�>=}Q�4I,��9�ʹ(�Do��pSvhU�/)��³!I s��g������0��i�0�+Ca]��}��Y�M�)V��ߩ�ҏB�%��|�����ɕR���/�;�J��5�!�Z�-���e�X�)5�3$�����q떖�F�2D>�|�XU�*�יU^O�������
�	j�Դ��yU:����~L�jO$^��N.n$|��AG��)�7A���&}����531�vWѾl�P��3r�yr�֯���pn�p �u�WC��n�!m�T�!1G�'�x�{D�@#�-!=v���d��%2��04�P �,�l�=ʎ�:�zu�+0c�����[���g�0��%^����?���f�5��Mè�e>�V��Dxq�,���KMRK��̺�"����RE"�e��@v����L�+]
�����+1H����`�>�"��he°�f���_�P�Er�T
o���f<v2?��Ep��u�H����l�i�ۂ-� M��0B����ϗ�jS3g�F�qj��D
mS�*WZ�1�L r�U�֮�%O9�D&�1�|�JEo�a̋-s+\�ܡ�x
�̷MT�iiC#o	����pS�H���w��&���l�(��-��Y[�3�  �c3pي`,�&#��h�p���6=�wu�ݟ�!~�x�rG|�,�CN������V$��$S.{e��V,@�VA�㢑��u�vs����,�'�2�Ɛ%fٗ|�	��}
�͐�x����߿�i����Ӗס_�U[]E�5��b��Y����M��D�Z�H(@�Q���+���/{m�E5+-!l�����{0�wsu%ڙ��5XV�꣥��b}89�3�
%��|~��,J���܏���Ȝ'J��.��K
�z:�����DS�o���d[J͔�� ��(L;J���L-�tR�7�!@z��c�oHwp��LwG[����R�`yyN`�i���_����ZQ��V�$f�t���Ǒx�aC�Y�f����I���BC��&R�܍��sc|;<���� &w{ _��
�(�+EJ!�[@�`�D0����ܮf�c��
@;M��o<v'dV�?�H(���pS����g�+T�	�kKT�3�ΑX	!TN81[�_��?a�y��M�e���)��7|�Hj�r�/�n����x��P��Q˷|Y+�ՆK�.������`L+�����I�#'ڮ�ǠR��g�v����_W~�:��Qd��#�\�J��J<�� 
�:��r9�r�]�ϓ�-�8�6*�&�7��>i�Wu!�u4�v��L����_��[Eh�>�����mܚ�M�;��,��I��W||ӀBS���p�p�[`�P��]s�����󯙸;�B
�_��k���1��?'T u��L���a�;NoDPH���3&?T�D�$�p�{�nK"MfZ��7W;F��M�lE3�ӻ��`)���dL��Z�,EW
�{ԑ]�fdF̆�չý�%lZ�R����F�-8�}+SҔ��K=�t��>U����l:�l��bm�]-�Ȇn�93}%dX��_w�Q� ����By�$4�t�2��8!2�4$�l��ަkp�K�6ٗ��R�S�%/1�T���x�� �$�'��rGY�֟m}s�*�2��lA��;��=�h ]��+pr�3g��#����K>��gCWK�^�3,3��r.*��r��D��� �E^�����W��N-�#Y�%"�/
�yL�[j��zq�F\��\��8 v`���z�6\�l���e6�/t��-�N��ZL,W��N=j9s��b�u��Hq�%��H���� �I��Z�&T���xK�ɓ9�_�e� �B�ĕSd��*�'~K��ɢk8<�q������y��ŷÂBNhF�|n�'��c$7t�_wTUy!��	"��G��?'��R��N����H)��'��mM@@��'���y��Z�)	<�_�E�)��������1l��`���>^~�9�
f�#ǿЙ�"b���b|Ϳ���������f]��U
�=�Uhڐ��H��;����HN~�No������v�ش7�q�&��,��'�D'���#j�Z~%)�p:{ 傅���րK���|��=f�E�Y�1KX��ucK�ɇ�1� vJޚr@a<���l����]%��
IXޫqI�v���U����ET��@e_`�)�D��~��	���E+9-�	�m�N�M��_TB�ˡM�w#��$�C�_(��VQm�Ot����z~ݪU����?�V���p���Ѱ&?捇[ �(~���<"����n֦Y���9�Ŝ� ��Z�x��=�9(��^��o�j�B�6�Z��7xn>J嵴��%���&�u�<v�����X��Wl�G�[��� �^�%��yI6�Ը���7�p��6&��i�jL�z�&.��9�)y�,�%m�	_��G���d6�U�V��[��"��L͓����%�~�7������e��)�Pv�^@0�@�E��0!�������[��woQ.�k���4E.���vl�IWc�^�\J�g>M9(��,88õ�3�tr����蕡SX��{u�N.�ni����Bl�)�gY.!q&ݝ���B�/yR��W��+�G�� ��j�wdO�'�;�.��q����@�N�-����K �-�W�iJ#s��q0���QD�.e��3hr�ke}riKPZJ#�ɨ-yT �D[ME��ęp����	$/) U���R�@ٶLWD�cu�Xx=�*�[V~���|�	���X�=�x����Sfr�)�탋=�י�'���V�ve2�WN��5�oŁ�$^JG�\��%lm�xֿ6�����gg�����{r!�35����%N�vX�P��
��0�b+����*�46�1Gx�"�b�s�	���c1�W1\�Z�vf�
��+�J�!�_3��[js�\��i�_�t�������˷2�6��A�B�����->n]�$��}��Y2�c�)S寽_یEHd�k���o�˫̹��؛��G�	X���0C�� ����S�a
*Aχ�����,��f�I��/��kbl��-�/�Z*EV}?چ��� �*T��=^�+ͭP[����.��|fX���+��9�'�����i�g�g�\l!�QG��r_���s�:ܡD���x4�'�(=���*"%Ɋ�Egk�Њ�����o���Z��S� ��/�y��+�;��ݣ�n ���I���CR�l^N��+��a,��:�h��5���'#�P1 H�[Z@�1]�8�@�H�<(q�*nsNڸ�\hE�t�������G��#��v!�9H�^����g�C#e�@Ej	��+��u���{S/c|�:#[�#}d��e�
(>�{:1���d�:�z8ҿxX������]�����Z���H7EB�xʂ#�@rHl��
rou2(bvl&�>��>�t"�r9z�h�h:^4���S�M!�7�N(vV9�4_��v�G�7+
���Z����b
ٕN�9������e��}��ƃ՗&F	��-;��3[ 1����Z�/&?Y�j�>��y�Ħ������5ߓ����N�RY���	� ����'��*�6��Q�����Q�o�P���EY_������.Q�a�7��/Oh� ����n<,��QJ�%q�jW~*6
���ҡ��S�ЖP�.�Hf�P�x*��! �p��b���f<����� �	~6���}��Wk�_�
��z�ף�ؕ���tA%���(�����W���eRuKN,�A	�żo����w@�/%���ps���F���6_�v'��8�k�rD�B����+�WV��Mg��K�+�Z��E`��Z~I��u�jre��n�3���	A,��ѾBˑjj!�^��dh�0��ԑ�p�|�HJ
TD�4�pФ�o��|)J��
��i���;g��j�!+<���YoQw�x�ykՖ/�cC�K*
��9��\�_<h��F#n������Ej3�:�� �>/K�
��!�*�;�gR���H]�+'�&��l�OM9�S^Ģ��<��|��~��ʑ�Cϧ���EԻ�Z~fZ��{bE@�"�n���eHׁN�Ԏ]��(�~�Nח�����J�����K��u�ʊ��M��C�ֈ֎}��4=�'�J1����+��bL��q�M
)�{GbBB*��:n3��\�MUu��%UA"�����zdܻ�je��U�Ԑ���������z>L�5�ym�u��,X����^T�:��r�:���Q��{ ,YiUm�l3߄�X�%EEi�|��I�^���?D,6+�qOº���f�ٜ�gՏPp!��⟣j��,��,�@͍�J�?����%�Sv#���T	a�y�O��:�*�Ҫ�'#�~���9���Vd�4̺â�7:�A��0NW�$�4C䧥��5Fmg%-�Fb6�oM�K�A���-�:�9sI�/�?�����dj+��E�&������V�А��p�5h�zf�s�L�4��2,`�ū�הym�&Q�1�;�b��{8�B�Hb�nM�<S��}	�.����mDO�?��~K�ё�(�u�,���~h�0�&�
1´c�pZ����PT�7ΫhV�T=�����	�	�}T�%��I�7^��˫�ls��q������޿��h$��$�p�w8G� �}6�t�t�+&[��:�l�lP�8!CvHP��)d��ZO?H,5�uh�]KV�����<���Ѝ�Y�L��*$���4��,��\+��y�Dla
m7�?��o�΀�[Sӛй/!���d:F�nb�N�H�Y�ĄdY��4��=���kک�i\^���#k�@O{�.;;�X��	��/]5� ,����4Q;�v��΁F�&\�8� )5Rm����ɯMy6ߎ�Ű/��i���LloZ�*��ޔ���ׇ�׽,^�sft*�7%]Q�!!o$83{��zt��ʢ�Et�����ƶ�C(�$��!�e����2&o:&�pD4C�*�4
�F��7��U'�%a:��%�(�3 ֙�I���fa��^�dr�?��.Mv��
Tꌽ	�&��P����m����ԟ7�"�BQ�j���s�.���B���M�H���s�o[�P���Md!S��eI��K���=`ٿ�Cyj���Y��>�6�B�L�U�@����,LP�*����$���䰦d�c�rs��n��ig� [M2�wb�|3\�m�8N��K�9�;q�fMxt�.zs��N����	�Q4�r6��z�$INE$\&�?.�\"�4���3��z��N
^m�S���y�^�~�$?�^8�E���x"f,`0�ͬ�gLŌ�����+�% �O��pFbh �}��x�w���jn$!L,)�\X��+��a�~�p�t��x�R����e�A��;���K=]��4jL�c!������,�\A`g��_�z��4|��й<�^��!�G!��yi�<=Ep�E������E��7�FL�L�w@�"��zW5f����ļ�fvr����# ]��Ym�Cp:��5w��G.�|�T��x�N��"�vd����g�1���"Z�@�)��cD�U�å:D����?���b��J�����er�P{ˀC)X ���M `D���<_���b���i+0�qnwO�e�K�֕��l�qX����E�׶w���'�c�g�[Cț�`����K+�	4la)A�kc��:�tzQVo�KXWY+k��ן�5>7�Q%U����b`T����Aی�ϗԮ	V�$ �)�cu�R�O�^���=�O P��Gh��WWiI1�i;Ls)���}�x�b�(�������	\��n� ���1�����D��_��2^$SI`7�iw��+3â� 9f��P�L���W���8~ļ�L��2&E3�	�#����r7�ҍh�@9/��!�	:�8���ݙ�T�����O�Ė�A-���9h�l��|�pw�l�=9t���,1���v��� X%Ok�
m�kk��s��qk����
.�C4�jך��Ʈ�u�O�K��us���$�=����6Y��Y2 ��+1�9]B�q��\Wf���)�ˍ��;���Mw_��AQ��N�[C�_4iS�r&Tt�PR�g\w�%Ƕ�hIvt{�__������hZ ���I��o���<�Z��O?���R�)�����M�	�^��/������h�O�f	����a�Jn!�A���,�~J�Kخ4{y�ײ��*�ä���"e�4n�{*�qh�Jĥ����,�C��l:}	8����6��8	%YK�7;� �f7Z���I�	�\Eb�<-qF���CMƎX�@Z�Yu�]�߯f��{�-���}B�p��d�mo��q���-L"D�)��֖��qП ꂑWJ�FdQU5 �6���o�����G�y�6Qan�E�[�: �H�#��P��Ϻ�h^��D9�/��^��@��Х�����P�*�FW��Jw�����ƃ��S� &GIc����S��Ǡ�����-���;��� �����N�ƃ�삗�/���dRD��w>�cYEg;��҅Ƨ����5��7�l\u�J����;+^L����+|Uz�r{Dx�SKװ9a�mau�Uoހ�pN	�rh.���m�/{)Db�rfG�Q� ��(�Va�J��AN��CcB�g�D�bgWe��<���(w��m��_&O�[���^{ ��棽*ܾ=#a�z�S�̇uj�\몕�F@�k���^��J?V$����
?�.��-g������6A��Ӗ�p�v�7�`�J|�ÅW�,ב�2�U�f��@K��E��������F�)n���S���2'����'�k�LAT���������G�����<'���[�hS�xu��d��ɸ�FuԐ��A:[zM��
��Q����);���S��Z�W�O�����*GLP��rk�i>�P
-C:�(h����(�Q$6'�=����=�\4��?t�z�ZJdc�\�Q���AY�F��� T��k�ե��kh8��uc��%5%���ԞP��ў�`}��P6�L,�k������ӍrlZ�X.h��E� �5rˬ*�\&^'d�hg[��>�"��axr��7-È�>�G��~���I�5�`-�A`�d�g��y����k����`��
c6�"�=qfԄ�񴕃$eI,���B���L걥4(��(/����u�Tw�ggQׄu=4~y[�3���]��B/Cl� Q�Z����@@��r��ѵi�(z��(o�[j:��G[����?�w�7�}(E���Zw�r� �	�/\a�@�.Ge{�bQ������ ʓ21�&�ө,_��6~*���B g��a�D^2���ݭN�<�E_�v�Fm����ݻ��0{ �����fRW;pb�Mvz�\�3�>��/��Q����idOGd�D>hg�i�i�Ѣ���N\7P�"-���N[o* &D�r�+����f]a�sS{Sj%7�J�_��H��8����)[�*�
�K�xP�[�����\V�����	Q�w�󹪬��3<���(���̳%|�>6!�����Q��6�L��`#�l�KA:F�VZUZ���/gA�-� Y��lD�fm�	ICJ��u��Y�?h� �&2z���b�������Im���x|4����L+ݐ��7�N�k�W�o��j���V4fN�Q�x]��kem��L-�2_u
�^�U���! S%M\Pm5��H�_��L_�� ����%zwvx����SP؊�ӡ�d�c.�"Z�U���`�,L�O;�7�ee�2�6�f/C_)������	��mkE�E��ک|���1�`$���Em�~S��L݀s��D��@�e;��b��Eb=�M�c� ������:���l��������4A�ӂ3}�@�����ff�9,�C#5�!���V�7ɝ)PP����р������b)�v����bwY�x�� d�^���wJ:������2c���{��������ϕc:�Lǉ! ��iR.������5%�!�n�d R�2H
:���*�I�Xm*�
5u����H��y�5j(
W�^Z9Oxi�ͪ�̈́n% ��%�����y��0�G�$�g^���=E瓮�1b��qEhW�-DT)/ }+�5-�z�+M�1ۧJ^�*q�����~/Kfb�%�_D�۠�_7��S�x��#k�9�5��6j6���s��Ub'n�l8�>�����Hr��ߜ�G�".# �����-2���ݔ)p3Ƒ����~��=�'(ܦ�����Z;@��'��C��7ڦv��K��wt톱��Ãk�Z!-��O��u��4�C�펝G�6�+��6�f��jr���C��qO �6��o5��E׭z���F�g�CiQ���FN8��_`�43Vu�X��B���~F���Q��R�jOō���6�c�1�%*&2���S���Iݍ���9��	�=B����wOӼ ��
�`O�����Y	�+9)q5|P�q�I�I�Y
���Ug"{e��n=��ǯQ` ��T$8�6���x��=�߻��2E�L�\(�虡��KLJ�"K���U5�'4�)���52[\9���¦�	�����W\D
��2Ck��Ɩ���\���8�����F���/�h�#��w!D����q{�k4?�S
�`_�g�I
�S/������@f��+/�<~;���w2	L�P�a'ͨ���g��"�bV��.��I�~2�/��L����X�m��9�&�"��CT�&�g�3k� *���B��I3�� �h~�,�a?�C�b-����#��+@w_)rV� ���:��p�����6���yc�ɷ�5�l�"���¡Ȝ}Gr����nFJI�{1�J���6�T8qN���_���ȶ���

 �XB�_�[�[㞑v	�me\^C���i�2�l�Hn��H!Z���s�)�?��?��j���.��gӢ��k�5{�Q�Ƃ�5�RϏ�>�q���Z�Ca��;*���9ˀ@g������o@��Fᄺʕ�q^�l <w����"�-%�hW�	�2�۲F�Q��l�����ܵ� ���~ҧ\��&�M3�gD�otJ�Ja6 �����^N�v�̠�����/��0{���FA�ә�6QW�Z���z	L'��������0d��kr�%�����mbnf}o�6���bɋ��AV7yکg ���������Q�w��n*�^���t@�0�t*Cg�6r�8W����i�EJ/��_ J���C�P�D�d�#��R򩕹� =!����7�h� �lioi��UB{Z�O�D��[ل�KPQa��������OA�7�R�呸�c���#��F�A5�j���?k�D���/�Sb'���Ȇ��1��:s\�5iR��cu�
�`L���,ӞW�[�j�
��nfca��4�(��H�ĝ����sk� ���Y��i��.m���k誧�]�t�픚���l��p!_e�3��.�u�G����m�n:�s�`'!c�ܸ�
��s�]瀔�	��^)y�`�W����o��֤����ǂQD�׮��|o����+���lJr_Ek��OիV�Jq�#[���L21�X��W+\[��B�nA$!t�u�{�����9㛕y52h3��@F':�W��J����R�pJ��B����O��ɼ�Vw�d{�]�ODh�x��a@�&�½�b�P�N�#�
jSj��|*\9�d��H��F�Ho4K��G_[��T���q��PO 2_��]y���S}�{�~�_�x�WX��N��]����^�x��je<0�rF,Q�q+�j����w���g���*	�����X,�tG>���*��5Ͱ�?Q�CmMc)St&?^�{��f4�� �=��w|ۨ)3�V��	�J�!�{�!C�� '�,��x�%�`�!$��pa�	Q�`��u�T~�}�n�oy�~ŘR��H�'�kj=K�k�#;��q�o�z�$E�"����v� �}�����u@���3Cld��7��LÛu$RF�����v ��̶02<a�42�e�w�"���3��a^� �F.���J���;H�.Z�ֈ5�����q��ܽDndo��y+��tf~��ٯ�P�B��CiK�%��bq�n߄�d�
d�`[/!��4ς��ʰ��˪sڿ+K' (X7�.�����GPĬ����9Z.S*���FnU��� �yy�lEa8Oh3z�NF���aXZ�l�\W�a gZt�2PQh�� �ڄ!.�6�q]X�B�u.ָf`�1�-]Y+���m��st�F?�QO�^�^^�}<~�#�xm��Y �H�<��R��à�!��PJhV�Ֆ59�����nȫ��c7}��MHNp��b���'���}�	|'�nx�u2�N����`�Ҳ�݀p��y ߮�;�PAd=*�⣢!�׭�r
',��=��r�t�(&7T�riK�؏s�cO 3�3z2����e�pq�N�4w=lT�z�� ^\��F:~0�{�����N��eZ���@�n��G��#���㥾�׎���=�E��"��<�2�p�tљX�r/C�ܳ`���lL����hqՏ�,��a�+Dp���	Z� ��������+x��ڨ���9����[�;���W��Y��3s����?ᷖk�����h��$����c~��]��(�=ֱss�1�-��Q��c���s���FpE�\R�����P�<8B���У<@���(5���i��J�w���bk�$�tv�(����c9A���M�n�_�_������GF|���Nb�=�J���;E�-��e(�&�1��\W��y�Q���X�:�xG	���������*~�E �S�KA��SQ�#�u�K�9���S������%p8��"cK�>��3E��ʈd0'e�VE�꠳�Jc���_F~�R��9�r1��a�6���\J�ď����� ����E�i�/�v�;��"?��6Q��\���Yoq�������x�r��W]?FO��̛�̿t��ג8_p
:�iu�BҐ[8S��58������-�_M��#B�6@�n�F����ܭ"���k��K�f��窰��
A� cm�Y �a�B�@q8X����ox&�� e��5<���T�G��0,�\�?k�D:��8�_t�cf#�	�����|h_?^:��CD<⩥ �����a(�ک�Y�tI�Rz;��"����;5��em����L�>?	�17�L����irb""j~C��\�-7˸��1tnI�&��F/�s[�#P��i�� ؔUP���g��A�����H�f��E���NA��8�#7��L��N t�s�������&�P[�;�B�)�&f!��\�� ��(����a���2_�X���$�����o��Wst��%�bn=w���ޕl�������(+�'�DH�>��,��o#C��[>�Ϳ�ȖĲh�%�Z�K�v��%F�LA�ą���Q��"�L������xɺ���
��E����3�>8��!���l���|v�?)���;n�`M�)_�bk�П��m�B�ç����l�fך���(S���C�a�+}5�7P{�a%":�����Ko;uO̗kfI��:���w���X��|��p���B]�n�O��\���P{�m(D��M$k|�_�p�׀ �\��KaR�Ï��J�5B]J�X��u��UD��*[�ڜA��}6.׻����gfj�����Sy��
_b+��\?��Qs��`N����}���xf�
N�����\��4h�z*�[:�P�z�ӱ�	���?��\f����mC��~9���*~�!����Ű��rc�����X�xAhI��!���]R�y>��n�xr^��1x�|���%���#�Z�o�d����A�~,�S.���-��8�����w�8��l ܑ��vh�1������=��f, ����R:*~�o۩��E�[�`��8�U��x�j{������e{�Մ�=�#�)�ǣ����u�	���#Jw�M�28��X�WT��w��𢽤��/\�~h-���@:H{�^f�ƃ��*bbq!^����Fs�ܟ���ւ�ˮ�PH2)x�^��K6,�yP�6r���1I���Pz�,i�G�c�}|> ��a������v����K~#w���Jc!{ �$���G^�~�J��IA�Uhi=�$����1�zv^��\�u\�c�á� @U�t"<~�=�l�.� "���:�L}*zh�K֏|�^7�Jl�<�`�װ��̐�ę�u^Zq�EO��^��h������og�T~V1�PKJX��t�QA©���_QF66 ����^�'v�RS�Bm\,���C1y*&�o�_��x_���3��Xन���ܧV�6�ϙ�i	jw��}��X������dE��F��k��UU� ���������<L���A�s�p��m�te1��(�C���>i��l�![g���s����:�g7���u~�Zh�#��%,�,*���*��"�u�jR�h$�z���)"�m٦�Ҡ���/��� ��?uF�d����Ǌ*�t��˛�5t7O�����
�T\;sU�~`��c�EW=u�s�8y�;-��\O��rd��s�z�����p��T���1���)*(��B<y��kk��e�� -�t�F�c�O,�G�a8�Od�XMT�h�kPm��s��u�^����&j��¥�X��m�F��vl�q����]'��.�o/:���x&�۩�Ѩ^iC�f_[���.v1U�v�XOu��Y'���d��
��؜k��l\���?'���<`��u" �O��)�+* ���9#�7���+�x���7B�����5���
�36纁o��N�W'Jߌ_�R)��M�sm�t���\yC\_#^�����C�r_��&������?�3/��a���<�������X�����*G��';mྐྵN�lB5�3�c����ws��U�����%���:ea$q\þه�S��������)�LT�;�/��$����`��S���j��ܑXl�Iå�0�>(i�g�ᬓV���:�.1�Ő��bM֋Ә^2�t�cy/�t@��=�f�;XRo�fk�C�{��Cp@ޟ}���ady:̈́�N�}{W�+��/�M����aί�B�o�����/:�$[��zI��@��g�@��M�x����*&X@Qv���Zv/�Jd��/���BqG�؃3��ŬUOk�{T4 lgw_�}U4#J���%��~v��;^j�����Tr{:�I��_�����q_ol�|���} �1i2kǐ>�Tr�V��n���`ۀ)ФOC�tt�s��.�Ïj����<����G� �vJJ�������A�m�p�k�ܐ~֞xh3�)����������C����'h�����P���S�-��ܚ���� P���N.I�ZY_�F��.0���;�@���XC4���"��zH�M�P��1H���c��=�P�;f�L������8�~��=u*����Iw|	�!*����i*�)��4�6��ǯ��Z�V{�M����m-6�k���k6��¨�#p�z�c��>��?�CeN�{:k0��o�vSafB�%M.������ N��V��ۉ������җ�`0$�X�@K��N���S_ٔ�?v)�EK�٘���:�i*EQ��w�]U���J;~����$������mR��I��w;�Sk���[O�X�V��/�!b ��$�/-|���%�*�~�����~7_�1���`�~�9��+*�9��2�.)R���==	bUdEk�E�ݔՐ�$�������,\&A�&�O�S�����Ř���%�M�A�r*��o�9K��LJ)jx���YX=��Z�ߓ����˳� �R������v,Ϩ��v&�_��������|қ�J<��\9�RC��[���U�ح�ޒH�#��q)R�b욷�����ƹ�ٮH��`!z��@߸p5f��wNdP~������zβ��v�+��F/�=;S��/'i�[�eet"�Ԡ�4�=*)cc���zܜ05B�8�6��o;:��[�"�;`n�"�0`tP{�tQ�j�W�<R�pvjT�
���e����l���p����J�⊄H��r1,�#�B��I�v��Zb�gQn��� ^�%��=
�X�L��S; :��K)�E+�.0�ڲ�;G�X�G��3BmU"W�4m����aS��?�;wl�"8:<#O��}���1�x��e�L7vI�^
�ǒ<(�V�萙��[9����lF��x��{;���7�Y�]/LYT.(ƚ��t|y��,<S�Nm8����B��&�8l'H.�J��鸚��0bU��̛���	��gGVA��?��+:���@�y?�~x*���\�h�	I��R����hy{�A/"RY�T��Ű��Ys��w��(�2zNHoj`���}��i�eK�H��;��eTEH\Q��),H�!߾I�]9D�wY>_kI�Q.D���i�7��vW��wXk�� �K3Fg�f@^t��ĳU��b�	��ȉ��z8B�`��m��cA3(��x+��\^��t������})��oY(ӧ�u�rx��_�����ĳX:�,�T]WȢΎC⚲��+z_0ѵ��/�ϵٷI�˨v�U]%PG��Rk^B���6w~D��Y)� �{�N��W�	���æ�֠�<��Z:����
L����b�p�}W�W C��!g��b)�&��s+��@���t��F�#�����GkX`cY<�/�"s���%/im��+�Jn�$��Q�ЕL���y&�1��&��ܿ�k��n�� -;|�(%q���y2�h�$� �&�Y>%�O=&����M���F��۷��ɡ��m�Iv���[=�r���d�op�s�X�e�F��"i2���O��F����2`l�X�܆���͆*Ͷ�nH�+\cV1�O9~�P|������ϐ��Y���]K��n�O�)��s�K�r[͸Ƌ��ѝ���+GU9Jپj���:�{e@)��V��(���?k�?�L ����5jС���׹4��$f�]e.�6�_�#^�ki�k$`\�}8C�6A�ج����w����*�����ߢ�;�-�u��;\g۟�Ւ�#���U+��j�*�U��Lv�D�<db� �S�oMp	�^�,��9��tnуם�8^��Lèm�k��J�4k���j�I���Z��໗ҦK�z��,�F\�l��"�S���<[(���s��0,Mg,�S+/~)��yy�C��*�6����_�s\����.�~��ӟ�(�^b`��
 ��Q��o�#ѯ��:;#,h�s-Ҧ)fa+9 ~�0��[Np�WsD�����Jlp?� ���EͶ ��D�t����	��aK?��^��Q��;r�T�N:���GM�6X�qW6Tngق��xb�v����i�w��1n?!E����MQ�I�+K��6Ed�}^�7�f<�I c3��9��g��B����T���*^kI�P<"�k�o&-b�ċףG<+*q8K��x�fi!�+bL�f��9���iŎ$v@�'ʦ�nÇF`��`��COk��l�`⇒��؛�,��������T��7���A�1#���&웪E�\hZ�	C�L�2�Pr��s?��5�"��S82�Y˪��['u�3k��������M��OZ�M;�o�c-��ͻ?~�5KsрԔ���lG&��wU�0����v��
�%��+�{��[�C3UNc�86N�c{}�W�$����3�U���)U�l?���lg'�6ȵta5̠�_��EX����+��wUd
�US��_�T�ChD��4̧IAװ��,JΡ�	٬p) 07ɯ�/��p��So���cV�8l8���Z��MZI�	^�l���g�6*����PQ����M���z����9#`�Ĳ�3� �0����i��{�GC��;�A'�g%�ΖԔ���W�<�)�I��ͧڄ���4��)�y�h'ĎM���ݛ�y��ӳ�t�թ޸�oF��5*��=Uܝ]x���8��p�屧Pg�N��l�
���-2Rb2����n-�1��W���;�il
���q��3;�Ӯ�a#�؝n�ܴy�2��.���4��U����BĨRR2&Y&�r�-*�˰2� CN6B`��
�9�}�1�� zqyȜP���3=��unb_~��tx�����+��6���@�i46$L�{�R.��=U)��=����ՏÒ߯�U����;5�f�f~�\.�@t�Yh�dP}�� ��I#�� ���ڞ��[c���q%���G���Ga\��Γ�Wx�L���~�VA�z��Y[<� }�q;�}��fTiJ��۠Sq ��Y���V}.�BW�|��w��\hsB�~L'W�|���Fa�d���H���L�@J^oƯ���a��-�S�q���pv�FfH՞��8O&��{H���^iY�[s޸}T�g؟�e[�z�]��{��p��k�6^�e�bE�=8P�H�&y��0��~�`D���1A����(3�E�3�����x�R�ȦAq��u 	����%f�K��]o�'�2��f��%I���B�lU�*�I���3�c7�r8v795���S�g���E�EOE���������dK@�-#�|F[E���7�`�t�%w���}�8�td1߲.mQ��F#�X/*�����l�I�"_Y����P��r�"¤��;��o,g�3,3�g�Ɨܡ3�e���4�;�o٤���E�ek:7E%i�����nK�'>�2�
/�i_ߎ�`5G����lM.�۳%��܃׵@�\Zc'�'6�Je����x�=S���h��Pɞ������81�e`�r��ʵ0H�^f�E�[����/�S��*ߖ��,`1��	��L�E.>Ϩ[�O��(�4b/�v5�Yh(��O%�ެ�R,�;V�n�Tӻ�]~~��2E���aE-��ȜN��
�c�n���=�USAL1�@���x�c�}a�:�n~���P�'i5v}����I3�U�����NI�s�zé"��=�H�>���5��a�-E3�������N�5�V��P�ΐ�Ѷ֢M�D*/L��f��k���c�_�FO:���"� He�A~�vʈs}��^�˧��qf���-;}R����9c-v��9)��R��hSا�\�N/��u�04��=E�?��	gң��z"�|�2>�ѵ'��Z�k*���~K[M��g�|!�Bν�cI����-{Z�4
AgB��r�u@O�ɽ�F��̳��]'���w:8v���<��� ���^�M�A:�S;'%��C�p6���_��#>ӽ�0�F�G�:C��Iܽt�n�S-|J�1�wp$9~�;�.���ۊ���_���
�ɭ��EL�?� U�C[��?d�Wg�:Iݓ)UIkS����qJ��.��$r��!
r�Mb���!0�h���%���d����.�$�đ��`o=o�Mߑ>%+C� O.$J�� jȜ��82H�ʙ:�;�T��Qs��JO�.��T�\�w�V�l�^
�M�v�[戽���c��E��	"Uv��/-���ǡ"�]́�Q���7��1+�d���9H/12n ��F15�g�^�%��)1w|�k���.ӈ�c��^F�V1�;�I��nh��KV�D=��j/�ǣ�����!�0���L���l��֐;�,���E]\���_��{L~��0�cH�E�Υ����c�<�n.g�گP��9�+{�P��U�T{�r?�8?��^�{)*����Q����o�	O6�M��y�B��iy�qY�?tR(��*Ě�O�h�������
p�Vk��w��]?�������P��WJk�n8[��Y+�M�����h�y�`��/؋4�P�\�!�ћD|�k�]�f����m�'�de���Gv����ݢ����Y�S��l��6��kG��\d�N��y40׫�E����H�,��:@�?�Ķ���'h��?�k��7w����\F-��o~;��4�3N�,��y����q4j+�V�:�t���¹=�xpt�����s�͸����E�*+{��|��|jsH���,�������$�u�ʼ"O�4�D�G�Uƭ��{��p���ܧ^�O�Nز ��%��w��A����ߴK����0q�1�F�mcm��J��3�/r�x	"F��M jw�)Avv�kz�j߅��7���s6ͱ}z.)i\�NC�\���@6��s�=	�A�FN�:˾,g�]ldZ0(�Θ�W�S�<����,{V�^n�GY�C��`yr��:��$�Ǘ^^tdRZ/�X�D/���G{�9!��ʙ5�,kh�$l�>ع����c�w(�9b�g4Ӑ�ou�� c3�'�K	$�^Lo��C%�8�fk�����~���6Jt�*@�p M\�l��$E���%V>�B5PD�V�)�A�U?«6A�Z�U���s7p���h��
���>#*�P��Z�a
S�����y���G�������
�]V���~a������?N�n�c��K���N3�b��\���v\�o}����ߧ �֠ƬıZC�` �x
c�" �7���(��f�Bttbɕ��[8σ"?�<���
�%M�iV�X�2����s�-16G���t���x�!�ms�Y"�Aw��p����>�l��m���=bU�Qv^��^�AT^C$	z�e��@�.Br�0�S��"O�y�T�҄V��XW���t��+�2����C��]�no	CF���0�Z�)| w��Q����H�}5��)��}^��T{J���.r����X+���&[�w�Rӝu��U�~���ݯ��R�"�h{7��HRg�j崔*1Ӈ�8h�r�I���O�:7(��<�.B���M0�������~��z�ػ��>��b#��� �m[+Za5��O��>���!"�9@{k<�:ٰb~є�
�)�b鎴�}�����֐pxJdDZ	�6!��\�v�u����kVJ��tS+P(AU�C(��]�K�!t�2��JS����8�_����V78�kbI�6���{�'sct�������}<$b3 z�)8mE�Y+��¾��TYDt���.���K�SĀM��� ��h�OL��t�T�K��^s5|�*
��v�P�}��2���pc����|�|�����1X����%��E����Z��l'��c�y6�lc]�.L��� �G�X�d�?�Ux9��	c��6~��fMPXˌ��F\뉚��g���@�a*�C`�69��-OH;i���``���HK�/�����C����!~NĢ�y~�B�:W�.+Ұ�n�c���+5Z��Vp"������%���|��!����{�
��B��JE䡕`�SN��NssZ�X�ku��a4��-cv���F�Z5��LK���"h�+�wLz�s�Ŋw�zj�c]�!$AE���N�l�/��K��e����s�����rfWi�o�	�~I(��W;@����`���H�����4�H��b�j��^�/���ꤷW�v$�Gg����1j��QZ��V��_pR�ȹҐ@�|R`��##yj.L�~B�Lht�NN����g����6rm��m��L�"5��׾����O��TSZ�j@�Bɶ��i� ��^RN��m5xeP�N�1����e< {�q� C��.
]I?F�����;Ջ�ƞH�����\��QS�OK���ݟ��^u��u˨IZ MJ�{2��6RD��+v�h��Be��,J�IZ��,B�� Am�D�?���a�ܤS'���Dޛ�$��B9��p���1ā����p�/����������'��k��xh���>��v{��m��-�!s$�f�@�bM�˛��gَBh��ypI^
;b#������J�嗨l�l�"�.�I~x�5q-x9��=Q/����v�$�6 �G^��O�c�bv�q�P�w5�	�������̛�U�lFB�K�zj��)�5	q�����f�R�Ey|�#i����,Be�RG*�m��G4!��lF^��+��;��7.�Ɋ�hXL�;'d0(�C�9��}sa4���1'�o�ţ�����2|���|��=�n���R3�YI�I�����x���fܞj]L�b��%ukWw��^N�=��ʧ����iX��~|h�j�m�׊�E�
�AI"N�J�h5r��-�7�I��`��#Uˣyg�Aہ��<�.l�K���I�	c0"�3����爒%+ ��N�b�3��/�yE�p����G��A���w!6�Wo��W�|��6�+��L1��]�QJ����
�nk�{�o��K�����n5����Л,�c�8�{<�$~�g��4��3ie���N�F�����&�p����Z���,<��ܮ�	�F?�� |���.>-�A5�p�P�����4>D�.)�-���p�R;��vځ[�ݰ����oIDƾ|8�w�m��4(LW��Nv�
��$�.lxH&�U*�LU:��I�avwR�h�Lk] ΀>���R��Ц�˲����##��P��T#V\'���H����Lg�� {2�]�c���N_�ʃ�C�G��4:�@ZÔ�h����	W�͓��^��+��6�83ȑ��������~�Z?���x�G�ҋ}ˮ�CI��m��)e��J��O�������GT�L/�)��L_]�Z���қ<�8뗋�G5`�����,%��x~s ��S���%��Uל�S`��.����x;[L1�ĸ��D����Tǥw�e`���R���q��ct'�T�,6%�S���c�p���{���y���_��?\sB�?,�z�D����S�6�%Oו�=�D����P-�A�$����/a9:S�y��'��+EҭN�R�G�=���8#IGe�H�Z�i��CP&`d>�n�ۦ��|yMi✡�*M�1b1�O����IrŔ3����`�5/'����YN|>�U�5��_���Wa^�Fy,�IQ$8`Yx��Ҝ�Ϙ�{Ә��/�]*����![;����K���T�l��-�}z�ƌ���ʩ����/�/g��n�3|l#X��'���*����6�ˌD�MG��������:�{*�a�A��o`�ƐÉ�m9e�Y�X�Nd-�%��K����7\�YQ�l
���I�hv����.�4�Ox�}9}9���ɡq�B �!�͡�3'~��1�������s��
����9��Xz�=�+"���o�z�HC�h�R�W��M�����'�*0�٩\*%��^�A3�B�=�t���D �Kr����S�.�	�%.�L"GB�$ƍ���Ÿ��@-*?V&b���� H�ڑ�9���ٛ��m�Qrh2�H[��>�5�?9��l��(z�R��D�:�	�`|M��j���'A12>�����*��ґ���!���'Bώl!�4O�˧���0�f1��d�}��
c9����@4X�0���"�at5�Q��g4M\�ؾ�J��=.���6b4��M;�Ӷ	^)� ]�vK�bd+ ]����%��:}/.�JU^گj�p��)&<K�	���E%k�� o'�]*��hrZÙ���x�4k���⩽3Y�jFKnu.i�,f�	����ç�{p����e1蟩���e��<�L\�xM�hF��.�z�:h��8z��i�lA�U�c ̈�|�~	�h%Ż��kR������*�9Ŵ@�@QctE���}���H5��r�X\���Z�]�2*�Y"��7�>�&�|�x2�S�2�j��Il�����p2{|T��<�7�x9ٔ�����k?W0�cl�"n]���:�t��5��MՇ10HzG�I�˪� z��T��B$!Ě�oT�N�r"OH�U6���bFPz�p�/N�!�n���!�no����}���e�sY�
[b]B�����TЀ6�|���U���0&=�;��C>$j^��Ք ��h����
8����N�|�T���e�E�_�Z�<]T��x{6��#(+��/@�Ls~�M�O�"�`l��i���#l��r*X���5�n�!s	�ec����Zt\j�J��xw�F��H�������=�(��[���E���C5|R����a+U�>�����\f����'v�{��'���E�:��S�^�x�N�.�GR�~�r��%%�w|h�,<~���Y�:��8Z��o�� J)Z�6\"�tt���I������ɵ�m��ӳ<�x�cBl�s��A�6BH,s��U�:�A:�+.��8Yӌ�@�US��<��t	�}7 R��d1Ñ����a�n�Tt* mȊT�voi�E/<��
�le��ϴ#΂@�I^e�L��U`�u>�s�|_e��+z	l5�])p h����o]�M�)K�ie��"���B�cVS�VW�;�����k��<r�k\zNh_���#.��r��(	���'����nB�y[|�לF�>n�U�}:�T�ug�	�Rl I40���X:��cF�J�#���A�K67BLf�"��K�M�]�5T�����]^�������Ŀ@��/����I�fVN1*Ɯ���n��e=�pR߾�f��t���;�C�x�V�}��p �W�[����V�#F1���T��*�/,��������HtU��y���cS�A�h5R'�F�V� �ԭ� �$��Aqп�:^�,Rd�qB���F�Q�ϼ�\P�&�HC)�+�'�+�1�o�����xJ[o�p�I�3^�m~�*
��#�\1�������p%�īB>���:q$���a��31�y=�𢙟�� �"�T`���kXns�j�� ���2d���Bߞ^NB�Ry
KV�H��uޙ`��3�Ķ��[`s]�]�dQ�Ʒ����V:Q��K��C��گ��w�o>tѪq��g򰹐�ay���	y�z�/ű�r�X��`]{�Z���ϰѷ���B�&�?�+��ڻ:O�'�:"�S��]Y?Mϣ�u7�7�1�8GV�Ţ�hK��i��b���u�-����7{��'�� ��gC 3�oP��(\&6$���'I�Ɂ�:~ێ�����1�������dA���ӝq��h���aI��/��t'q��r���Ay���ɡ�Ouډ!�3�,D4G,�d���O�qa�V��|$��-���=���y*�^�@�w�Ƚ��a�L|��I�=T��/u@?��g�!2��b�~A(aE�1���<Jǜx��z�S �Ya��@�N�Z-�U�6�pw9�֣����5D�1�烖3ף<�R��}2�3�-?�L㭗U���5�)�y���U�Nw��;"�G�UG���h�����$�Lc"!�5�F`ɾ/f>��_��`
?�%�����r�t
�.�)6�$��ֻ�7Z����$9|^��)�Gߚl�����w1rA^�TYqh��b�=`{?>�k�|b�������RV�)����d��o@�T�-�� Xtm�P���r��&�!F��4$���Q;�����4bi\-�s μ�UJ�yDX���
��0���u�ft�߯uqMX�s�:����_�Yg���S֡�k+��t��-2�{h�J%=�pg�Vs^*��%��d� mG�;�ʛ�8���Ysj�M�?ݟ^^�w�S	�(���B,ʣ��e}�����MO�K)���-�߁[&0�wAȘʃC�8;7:TAC��$��SP<��4�j��-��x��i�IE�h� ��n�k#=��o�9S���/���W�m��RNgP�$��1��'��-�����ic>s,b����i|�~Ay$��)�ND5;�=��&����_��Q�/� ��6�w�;��I^�o���z<��}Yzk'I��BH��S��xZ�@�,�4�%9i���k&��)d�Uv@���m���LJz�S��TJfM{Um��c���oc�Q�'�́��d�[����h�k~r�9�*}O�B(�+�m�R���b@d�%�gn�S��Ɨ ݟE"��5�؊����(�1�@B;HK��1������~�?]T�I�� �"0*2�G�I�m�a��,���ݕ�[�'S��*��kB�?Eѱ�U�E����UTOjӕ̲���z��BQn8�4��5�$�B<���?0��(�\͚{}�c��Թm��F+�u_��Mdk�P���:tC��h�qA��s�}кl�8􇈮��/��R{�ܺ�R��}8�f|V����.QΛ<^�:��i�TƠ���^|�d&�1���N����7@9�G���&I�x�,^�4[.[��$<�z���.lcv�j�.�*�7�1K��j��]B�����\V��|TQ3m)��W��u��A!�nS�ǣ����m�B��ޙƍ0U��M��)d!1��V� 2 ��,W��i���9��]�h�������=�^�6�d�1O��ZrT.BL�cs��9#���n�7&d�4���Հ��R�i��N�J�we� L �}��m.���Ҳ3����0�[�Q���O���,���x�g���s����W�d��t���<��W�TJ*A�(�8�nE�h=`)y&㬠 ��]�g�Gԛ�Q�FX�Y���T֩�A����xF�I��?i��҇�;�g�2�
P����^���n}�}vCK��Xc��d#(Fz����;�+�����b��q����uY���p�E���I�����1:)�oZ���Ќ�V������ˤ[\I�\M}��9�PV��Z0�j&M�2��`>�#ǯ���Bh���~� �����KE�%M�C����@��}N�'�K!�Z�cpytS-�6_l=e�����=>
�}#�o���E��K�Y[� 	�\3�{�T����'Ls"�)���JLإ.��9��?�Qm���@Y�a:m������9"\����G7��d?�~���f�$�����^%�"PF�%}\��5%P�ӎ*��F���]�0�P�#&����G�۱�G-��+Ҵ`l�,G�<$͜� �2/ŝ'�M^
���M+���H�YCG�f^���~��r�8�4tB[�Ɇ\��ڹ1X���!��Qu
Od�'\hx���%�d��IF�R�!� �~wP���DķDow�pZ*K���C�,e\�-���T5����`��9�]�-��_�@��#�QI��"5�b��	�X7���HC5�b��֊��ʤ��E�dr�`?�0��˴�O��
��pȉ@SHQ�E�;'RD&
�.��&+���(:i�/�aOaZ	oa�5��4��o2��0L؁��V#�,neh����}M�K
D�։�cֺ�TX G�"Hp.�sM]B-�#>M�� �m��M��Зs���R�سɱ�O.�=�Z-�CD;���NV�B�h�q(��0�lYi�Ҥ2FY4�Mݧ��m��9�f��,ܸ�O��S��Ҝ!c�~�t���(�f�����-b��ëy�^*�1k��Ox�&�Jކ�"J���K$LW����o-.5lM��/z�_p�F;���;��0�d�0���{Z�eY�ɋ���.�N��P�<m�#Pt,�s���V`��>�֑��v�E[�[E.���B����9�a��j�:�`[��d
���Q�)���k�k���e V��5b�ܺ��1���/�Z�����g��w�i�5,�3��IOa/"���
p���:��<��+	zRAD�X!�3��+pw6��)��a>�<�{���)R��c�:sU�H56��7w��6<�����i ��z�s��0tz�"�D�"�j�sl�l{�?�D�h��[r8�_p�m�f�uǟsֲ1~�@��B:�Ԁ6zj��Ģi��&bT�J2 �(�����V1���ԟB�z�&"��8��D.��aO��/X�8���
KJG������u��Yy�����)�x\�c�Kkj&�C�z﬘��fn�"�Y
��w�,}�����ƌX+'��r�}�lѼ���)����8L��x�f����Sw&�܇�����@�o��U�-f#�7N��t�P���N�y�5C&����M1ߏG���<�*��<�=� p�1^�9������J+��sc�
��n� #�/h��ddqO5ʨ����6�9�ȇ�(�k�1w�ƹ)�Mh��=��=X9�w�"w�x`����x[(��W��]7i7=����B3���zo�Х������j� ���	 e���­�>=��i#��!�Mf�2нtLE��9>�r�촷I3��2g��Q�p)C����ϲh�@H;�+�.�yrY�:�cT��i�^�i0��[B��+}��c_L��j罸m����4z�!���+3�M��;Τ藽:4Ub���NODT�����|�sJ�����w��rT��Qz�SS�?��S�K�E�WǗ���X)�B�hc�KeN]���*��@�:<��L e�`<��U���L��@V|k���_�l�Mxཻ��W��3�E��*�1ۧ��/m�Kp��5��o�a�/w�<�x�B&ɟTԮ,��q)�H6�{�}����[C�
�;+��Yݚ�<�;4��'��V�G������b;$��t��>H��� 5M�uL'����%���M�7���bwu�c�}���ɋ�K��ф����%�u�O�H,ϺW?k8ǉ{%g��A�������`�d���ܷ����{ҖE0�{�
�
�SK�	�K[1*wꙻz�Y,[�S��rTK]oS��U&��t�H:��-<�?GT��D�U�d8�
ĺ���&9���V*3R���Gu�ێ�#�a�R�T�n��60��ۖ�q��& �iN�rv���qѸ�T�{��I� v���E|�����˜�E��fX%=�n�h�k�Ծq �����iکt������S��SB �K���¯-<�����R%�K-�������|%��.��C���+��ESf�q[��$ϭJU镑F����l ��1xIܐ�-��\:`Nk�z!�b�keܵf�l�8���/�S��!i�Xpk��>cJi.4��8����B���7�ɑ�#��b��.�QX���H�2�0��w̪�@֎��/]����� ��1έ<媽{�����5��4�bO�6۳�s饦�C���M��U ��>W��I|%Vӡe"PNXB�n��EqR5�ٓ@�$��� #��dۭtie�P�XٿV��lg8�A��������l��L[ԏ1�չ�z�&�FT�!@�B�q��bi[������B|�M�M��ņ;d�.��?��[.����?�������5�����'���#7��Zo�@H�7W�"[o�)���8��S���.�	E�9_o�i�пF3ZBH(�~��cR�*i4I��]}���纨v"yͬ����3���P�xE!���ocX���V���>�r��O>��7�^|$O;\�	��������G�w�{�t�~$]S���j�x; ���-C]S[j�����#������K������ ��=�Ҩ3m>�*�ܲ]�(f��h�v&�#�K�]X���b�Ke�Z%�<�lPrn�w�0�n
��jD�)�$�@�,����"-qU�&v&���E���9��I�������
��3��ݽF�ڥ��^��Q���_�Uc��zR��R@�sn| y���K�F3T��3Dd�fv���(	��P����V����"1�v�U�^n7O-�2��{�-�U�V��������`k�c�n!�0�������6��l��o�t���p����|p�tJitl��ף��[D��oX���v���F�t�6���dIY�M �'���$%m��p��`�[v�fx*4[B���h����aǼ���������zdK���EOi��Q�mR���r��v�-�@#}5o�ٯD��O�qU�� b���XX�LS��b����$E����~��$r�*	������Ẇ=��Z���w���m�����1��0�>��6�Ѹ��LȌ�e7�(�}�~���@1{	m|W#�!j�����Վ��C��qè�Z�#D���^z���sk���^�ԃ��c3�.+0����(�S�B:G\}�{G��ŉ�h��n��⼏e��U��D�'U7)�0��d��|��^HX�A�	f�Z�հ�� ��p+@�
�A�cp������d�����1'��LS���g�%��-�x(��~��g$���mn����K2 	�(2|2��y����nIC��a��ퟞ�*.+sC�j���10�&��C�˫/G�F���0�j�$�h��RЃ}&������rHz�<$5���\���~l��ց+���Cx���
*��FyBov�
 ��q�}Nv(�L㪒���F����a6�="�)	�����.|���sg��z�
����2	j��!8���X��΁UΕ�]��}�T-��Z�F�0����p��M�4�a�k���Q�	�P���9y��"�0P��1o�>��Cm�x^�J+��(��O��P'����U��xDr�}��*��܆����(i�y�	kK]��0�6<�A"��q���T�]����6��M��{���^%Z�@r�lZ�xH[�n��R�Ek�-UH��yU��/]�C�up�����Ïpȓ���H׺�6P����'<�h&�d�~�OP}��ޟ'�{��f\]�	����]�v8�+��>�w�}c��p?��)y����Z󓔏y#c�� Q�H���	r��zf��O^q�wܩ�ZLqm9�X c7ʆ��L|g���
��&��δ2��Q�du��6��ɫc�}@Ό1Ϗ�.'T�x��_�h1��1ſ6�z��*��_����x��.�ت��t|f(��g(���G��0������D��?���^�I�r)�k���oW��X�ɴwyshۆ��d4�����'����<�ل?�+[*t�u#gW��6b�`/GE.~}� �MFi6�cq��Jn`�l��3^ǽ��?$X���w�hR<U:HL�t)�5/��-y�Z��v�A-+�慍]��U C�F���b��}s��G�0!]Gi������B����q�e�� 2Pu��,���{�p o�	������S�a���Y��<�:�/)����j �z��%�y�ih�ڿ����t�n�$�3�@���'I<49�ۦ)��o<�y�5���iƁ s�B=��yx�	��Y�l�B�d��,0�1��w��J����v�^kg�~��>���E�6���N��ظ�W
3��kK�{,�F�eU�p/l��� g�贬v\D�C�@p]K����G!V����xS�M�l�*d )'cy��Փ=L�Y�C�x9L|��cxhc�Ϥ/��&�nI��׆��>Dſ%X|�:&U��d�?��F��K��}�����b��f˦���˰�	Q�8ƕ�W�b�k�̵��`��d�
������DqJ?h�0ھ/E�J��GW��O���o�
&:�V�f�Cݺ�*LO�,�}Oy�dh�a��h���B�zp��ɧU�ks��d�3��#ͭux/��Qc�U��n�ʚ_�%|���\^�G�3X�(�P,�i��f?�`@���5*���2	�D��r��s�"
���_܃�aT���yԷC��%+��|j�	�PF��������$��xu>�sTE���8�7���c��S)@�O�O�y�����+�?��!jy��!Ӱ�ז������˔ڭ��E��|��cSW�t�"�\j����PX����<���!�M�=�� ���/Sq��jr��3��$v��6]����SbV*6��.pK��F�����&�ȳK����RU$��8�������Z�g{ڑ�hg_��-$w��ڪ�}���"3����?���GV��|�8�r�l��e�Q=�����q���z��C��0\ '7;��n&��C~��Y�y��
�[cM1Ob�������YG��ꗞ�/������Q6�}5��]�f-ƿ��#�4Ǭ��ʖ������T�1۔��Mt���.h�к�*8�9֎;�Ҏ���E߫��̯<aZ�B��"�y���wq�Ek�C0�{(����]�|���t���F�m� 9���P+1���j�9���W	��|H�yAJ:Z��3�B�d�y��Q�s$����+$&M'��7�:O6���ӌ���2�YT,M%X`9СOFU�H�����]ӎ\w�T�� [�P
��ٺsXF��o�*�RX�0����&<y�	��C{���F5��"�OMg]�B+�ϔD&��p���/�7*%�A�'�AtQ����h�ru��j[���vKS�B��	�hL��j�?0!���"���Y:��8Q�FQ"��Ź�(����ᗕv��C�Q�*�x�E�Y��R�dZ�w>T�i�������F\�)�UI����1��Nٛ�����_�@����M�X��H��M'#r7��JE0\�^�E|�uv�zH�+�䋚������6�,�n�E=�-��6L�E/&�`���b9���j�w���.�FK�3Je³@O-�)���D�s8,(���'.a�Cg�R�.��������u��[0�Ap>5.��
o+ɿ�`A������;!�E (�VY[n�|�	��h28���"��KȺ|9@N�����"���!�:.� �&<G; qs)�@�^�iB�w��+l�%�]I��C["�g.eu���1�آ�T?ׯt�Qq��f��aލ�d
�R�iafBZC�{`5��b��".�M�O���Wf�¬�f�90�I@e�*|���	��B�x#�G��5���U�&�BFs�I�/4�"�5٢4�`:a�t`!�MW�l��i��򿮁�y� o�)F��?�ٿ�y���M�HN����j�W2��R�H��c�S� 8�I�@5�;�����jるG��{4�:-�i;ί�e6���e�V)�,I�!٨q�2�y1ӱ��-�S�d������Pg�DN����K����7!��ad��$s9��i�������/�= 8�+Vq�m�N�3��8���q�FLt�*�=��E���v�[=�a���P�c3�D�[�/y��Anhh��K�g����!@�9S�i���!Y׿����*^y��92�jh��k6��]F��Z�����m�m �G�a	hpSJO>VQGT-3OSft�Dr��e,,Z�gDy�@��5�?OA���q�&��������{Q0�r /�R�RS��c`7���J��9[h���U���9#�ՙe�� \NlUT ��ꔨ�JG'������S��̴S_؃g� ��^O���a�����ڱ�ΏQjG�;�V���IhS7�a�;��v�h'����s����/�.�{�������=����7AK��Mk�`��d�|i��F>�����0�?������Pz*���x�$KLS�H����S��9�<כ'�v�h�qoX�,�����#��������XT��'.�~E� �*g�Qy�i^۷��.�.�HT���1Z����R-��Y=:�'b�qh�����v8+B�%�/B��9V�(ܒ꫏ca��jƮ����d�T�T�VA9<��%�7m�|�im�2p6J�G�B����9	U+|��S	�񬠟/3�s��s�L5����r��n%Xe�'�0��xE"p��d���?��|(t���(�nS���o�G�URn� 8� R"D�vp�C[iL�J��"VL%i��e8m<�����"���Ԫ��
D/;aQv:
���_�G�ӂ�M�`��/�&/�^X�Ӿ����� (�yT�c�a�����_[�r�|G"`����Q��~��K�oє%�vB��N��b~�6��Am�3��0���Hw,p� H��^�EJ�=�S1����9���ـ�ȁ�����Ǽ�eIQ�0��m���Ɯп'�3��b6�pU�C���rfp��d^^/%�R���ԵJ���b�x4�����j0&3���iق�ߐ�t�6XݴC�,�x>Hf��f��b�Du21����6a��ҩ��f����_��M'�6�U+$emV;Xt���Q�Yze��C�Cf2H�b���1�O��J��R���h���!CL4��P������A3pX��_%�Gb�D�幩���X+9���W{�����o�J�i��FZF�	�#[N�mC��^�ct��0i� )%=��3�h|dv�Sؠ�����	�-Z�6��J���>��M�r6���������X䙍�������J�8�luC�������G�Ogݑ��C;ߔ���.nY;"���.��g5��吆,K�|nW�Ou?Ul(�N�9Y���ꂤ�6���U�2ȡ6��Y^D�s�w�q0���7���zv���w+}ԶgFm�U�c%����(�Qs@���d K`ٱ�(�s�=�5�4��U�Ɩ���:��l?�R��B�-"���	���m�d����.�­����)���L�W-��M���QT�<�*�<I���v�3ŕPO9z�ew�E�1�8��Nh���ș��k(^�=ep6G��/S�w�|kH4�����b<�����?m����2�C��'���<L�ln��$��lw��(��Ҥ/��I�h�`���6}F����e�:fv�$1����#���Zˆ	���i�yƈ/�&D�)�;���
��(f�:Ǉp�\������y����H�4�5ʸ=X�����2}Cn-?���$�����{Ʝ���i�ޕ�d��̸�<�� _R�P�;���Oy�P,�c�n�� ��}�tl����G_������8��h�̣P#B;��(;@!�RD>!>��mUp�*Jυ��!�����A8��Iv"��h"׫9E��<M>���eŪ����_S������k�� �)%�y~ڴ0�+9��iR��H�Ng)t��:�ۮ���K�������L�L�'s˒hq��D�_��p�ş�7��&
!)!p��R�����-�W��&�������Zf}�9�-�9N/�A�j[��ߢ�T����>��IGsv�#��Fd�D�=��?�Ļ���,nCE�2h�y>Ê7]+�q��+��ʖ-J#:��B�Bc݄&�*�=���+=��I�4X��hY�b6��#�J�f���&�o�-�� ��7������ɧ��Wy0l5�<rKH����DR��+��4fvܙr0�F��ǎ��)�cn�k.���^��G{$��6����ﳏVs���f�p���%�,h��N���P�A���O��%6�gm��w��Q�����a�0�0L߻�*��Oj=< ����0(F�����z4�TP�����V��Z4�!"%��F`�HG�!�8f*b���G��6��}�^�j�]�x��4�-!���0��Q"N���H��t��؊L��v��z
�u��ȿH�{	�<�N��w��������%�/xsȱi�����Js��~���DfR��S%I�" �)��a⊖����Q!��W�z�^ږ��3+�"�� ɯ�㶾��~��=���Χ��)��ĵ������y,G���ȝ(��CmUc2J#"�Z���O���2h0h�4:e��53�Mu���n��K���L�{m)ר&����b:�+��i�.@!k�'�p_O?8��ɍ�Ut0gR����F���Uq��H%%���-�n�9�\!�3DIW*y,ݴM�e��ۺ$����x�	!ŊezL�߈S��ړ�duPw�ꦤxr��	o&^��r6��Z�挣���-]���M�6G�W}��2Bd��K��k�i�&����Oj��n��:���[�߼j��ӄ�v0��	�l�cZ�}��;8E/l��h�{��a��� 颶�R�*]>:��E� ���v�^�.3]��V��߻�P*��m�r(P�ޞ0�}*�3����T?�p�Q�d�����S�}�����z-�6�h�OAv.������3.2cq4�����.c��a�ç�Gpo��G�;� �.�G�,��2�oz�2N���@u�����C�K���%�Q�Ps'Yz�G���9���9_5����ެ�'�=���j����D�#�(��s0
�` ��dY񍪃q{��)�W!��+ m�d�#��9,")�.�!��|9g ����;��d�I=JIӐ�*��t�ʱ8DB"�+��FZo�ɼ�>��<�:��#�)`B����w��b����	�'Q:��"x](8��F�!+I�D"��a�,�mS0O�>����;�ۂ�u��H+qSD��ښb�igqb�'�~�a��#���Ή��U�O	�#A�}���c��Ǐ4ݣ�(L�p��֫��۰Ĳ�:��t�;5��Ҳ��0hPۦ��|j=}�����/ ���QS ��%y�8vT�)ܞ�Ց��79g�i�� ��XuU��-����8���HRY9o��B�EzI�_�<�B���w���y˝���R���#�s��i�
c�!oI�oN����z�)�Ţ�;ќ��링��:�/��j4X���m��C���&�d��Kލ+\��.h�it�β�<��vf�&{���Ǹ{/b�&ch�`�_�7]1[;mG��aWs�+}�p��<�$u����/J&f�`��d���tsQp�cw���޼�l�U���6x��e	܀�τ�	z�L���U����a*�����P
�dE*?�0	�lc�Bs,��Zg!`�#�5���[	�~�-����4���M�Ǹ����ṙ+07 ����\�y<�e�qy�R&݌K��Ej�Ҟ��n�_-c��L��	>��,�^�b#?U�31-���Ǭ;���O08���[�@a)O�?�u��������u�9�6�
�'����֜LG��Mgp�-����_\�����q�|��0��7uU�w�II���n|Z�q��>�|J5y����p��K�Q�+�R�GR�v|�c�6�OB򨠈��447��������"]
�q�.�Df⚝�㮩��W�눶G�B��m�zTe�j��q+�  �!/%��E�
g;oY˱��f�Xc��4�g�c*�r����&�6��mK�4&O~�o����HY)�Z�|#���~�7]ۺ��Dѯ�����G)��֦R N����"�e���?��?;���f#ʒ�8��ؘ�ȟ�a�еjco��r~JD�|g8��nT8��2mh�Qҁ¬�ǝy�9�A�}�|%��l�j�'%x��P�B�*�~ߝdx���Qm�o)�W�ba}m퐂��߂�c0�l	�9U�H������R�A�����M��m��<�i[�wl�fy���_�ܨ�[Б%'^~O,'��S�7l����pwm��:�(�c�� �,�Q�_D�eO5w�L0%�ո��y|�vE)H�7��J���6���U�@:$�M��]ώx����"]��}6�U�B���	a�Z!z.,"�U'5v����ы^������r�\;u�ф�u��l(o��	�f���}�>Ys���_�E��K���*K��>����*������F��G�t�8�UN����X��TO}�DS��>4ۧ�v,�Q�o��H��w��/�w�:��Ix�o�o���1�A�� ����'q[��B'`"��pj(J.�I�L����e�v]SK�l�I0�8��Ԉ��>����]v�G�ew���T�����l��y��s�,wz�M�ߌ�ǦK��N�����W�Zd���ZTz����G����3-�э��@��[��+�X���ݏ��y:�]a}�<3�� =�t#r.t�]dp��r�uj��-BZ)ȿV�`�ŰN=��-,aE�Gu�/y�i���&���w���K�U�������
�g��P��+�4a8F�@����o�wG���8M$v�OW���n���p��wF�H:f�#"�d+�
y�#�x ��z��l�R�١�k��ԝ���۵�w(	aT�n��\癹��w���˂�JE�����y�唄�	{�c&��V�)0�0o�ɽϢ��X���r����`v��xV�]�a�fj�Pf*#ԥ������s�\���J���9�f���.X�F^B�@��f��{�j��U{��T`8zԤƑ��^`�q4���+*��`p@�*��+�1jZs�l֎�O �12�pJ�=j��9o<�͠j���K�T��MQ [&���	K�nq��AE�b=%y�A���
+ZI����e�E��V���b����`�&��F�aY6L��U����S1�P$������w���׏(R��N������oD��M�p�^/�)��^�'�<J���.�Q��GOdZ����m��s�h��): %���5@:�3��8�4���x��=I��6��M��H4���,]6��RF��(d�xz_�VTua��U2,q�\'�e���?�&(%��̾��&�@�����ls�^~'��a1���{(4K�b�b����1_E��I�Y�ւ�&~��yk�GO�n�dtݗ��i�ׅ!�S�Ѹ��3W$��)�7�^?����~�r8���n�7�u��;,%㋤���W����/��H��,F+at�W(��m�7���
�f�9d�4�G4U�%Z��w�'�R�څ:Ъ�4@�<  ��L2	�����Y�"vPnr����̔������\�&���"S�����)c�����T]���l�՜#��z|ť�B���h �Y���C��\������/�Ś|_Q3<�T�k����  ����%�S��A�g�+NmT(�Ɨu�mZU4s���WO�*p0K�ӯ���o��"3&.��8>xa0���V��HXZ�+�:���%^Q����	Y�~3�b*E@V����z�.���M4�D���X�Q��Ǜu�q����	�@��S���@1��J�A�3_q�#
�kş�j��X[kh�����wK����)��ZZ�!oc)�mJ���h�P��5�e��'d}-��f1�������~]4/�Ŧ�5Vl����Z�F��AO���0�^]1)DE�nD���5�s�!�zB��7d��m�{�.�5���Tz����t�rP��Z}�Hݨ�ϛ�7��P|��A 3ooni���"H�s;;����e��U2��뾵�jp��6B4����3��sG�*�e8a[��R2�?�t�X.�
����`�G"tzޱ������S��g��՟�1�������
���>�n�L���Z�4�3w�>ӛ<� i�:��s�����$f;�.��c�$-Z[�CF���x�O����}��3�rF�A�mG��
,��{�W��"���ǹ�H��{��5��8�-�,�����<��D�V<�RGY$��*s��@t-�U���w1��J��f*�OH������ފ�eR^��3>w��	{�F���u�ڕ�f�Ne�t���`\HbM���R��S��|@�S��pv	����t�5�x�����'\C4$����q%U�NT��p=��~|ca;=Ȑ̔��n#t���cX�}4�=����C����OH��`e�!��r��W� ���4Y�E�o}#�ب���J uG�%(}T=3��3�<l� �R�A?G�Cit~����sG����#�~���F���B�'�r�L�>.p��a��钞ܙ��B�
���?���u�<#5dF���.v	>\ǞW��1���V݁mC��Ⱥ���!��UK��ǆg���q^m*yl�رECԪ��է��%K�XrN�� �N�_��N�2s�[?Y�xzq���kp�H��v��"ա�CFD���t��9�����Y�N�8F�^��ꢉڶ=,@آO�پ�`1�����ra(
�q�q�31��5�x��73N̒;̇H�(�3�%q��ڰ"�[#����P	g�S�n�8�Q+�3�P̬��+%����ͷOE�B�̕��*��Ğ/y" ^R8��OĞ
!n,�eH�(�ŽnuAf����� b��!p�1���5����`^���ϴw��w{���"�I[wnx�e����~A�ǥ�)��SHW,��z�(�� im~ٟ�RV�P��ւ;�ӎ��I�p7��]�K�n���_~y��y��hp������]��M��U�o�G~L��>�=�}{�<�ݕ��~jrH>T���"_��%AѼ�{�8��f��]T�ڙ�!�˧-U!ҰSR?l�wN������ԶZ�� ��b����
���^U�;�yT��L=#�@�l�e��Hh82 ��Ba�C�2Ζ!�*���}��Ѧ�t��=u�G��+�
�W��sY�]�Z�R��[�S��?��:�u�M5�*���Ỹ�$�UT�TCVZ�j��i��w��E��T� ��p(F��E]�vM,����)��[��Q���-7m�%zg� �j��@��Ea�/�V%rP��L��zrnv�r(t_��gVB�:���Z8� m��VI,�r4���s��(��O)�cz1��P��T�	ɻH�!N��3�e�~�J5�:׎L�n~P�3��;��z�y5񱹡�S�/���ʸ�|�[NO^���-�Oe�V�WH+*���,�����{�8T{�Y������m<��$%�j������^���J����,�j�kB$����Y1R^
�+¬��-����.!W�r��$UI��á����4������X{ռ�(0��'��|/���ʦ�S�6�����]�?�󈉿*��?ImÒ��1��/�*�G��Eo�$�S�kBH����ɦ1�����e��Sx�m�a�P��J��-*��^7*�9c�Zb��0�@;�Ɨ'@�޺IX���I�������&��ڦ�S��^�s�~T' � a3����6P���"�����X���C�coI̺L��>DYb�7r��N�&�١#Z<?���4��h�N��ϲ��-�F	�N?c[`���RH��K��I3�;���2:��_9	���xeT��j)9#g�<'��mmQ�#�ERN��qTeih���Y��wG�
�'�?�ƳA^*�kt`p���zi^�����$u�3	X�ڪ�*J=x�v���P4vጱQ����t������n�"�rÐ�y���	��tգ�zs;/e�;`��FP����(%	{�bn�U�i�	��[OuPM��^�XD7�v�܍f�yv����0϶H�������U7s�/w;C�Oۥ5���c��g\1`АH7Q��RͲp��`cքϟ��0Y�kdER���7vC"(\c��!�Wt� ���X�|�<�8b���Q��9�ˋe�T��]r$7���ԧ(�f�-�����X��&�L&�=�"ebh�� ��_-�"|��}���w�]>t4�$���m����7:���f��R�M��O��5Iu��"��>?���Ե����l�@�J���D\Ə�Xvʅ��n�s��hD�(�� m����P��Tk\�W:G� ��+�sמPe��$���f��e6�r`q�,d�ڿ�E`�/�@�"(�@X���pm�o�ެ�g<�d5�s��6���Ci�c��a
2����(�htZ�d��bZkL�Yg3����󛧑jfC>L�4h|��K��Ϋ8��-��=:��^��Î�׋�rmq�:�F#�\T�.���@joc�4��yo�~�)ߩ1\u�ֹ%0��^�L���E�}�$�h��%�_��0\+~���#5jN��Oc�@A!4�|��~(ő���YNb��3���W��t�1��!��~���j�O<:�jqCK�nDU�A�v�u�ou�J��TC�_^vL�����9�=y":V'e��I��M1fl.��Ԉ2���L�!΁�M����9�Arx��F递m�m�Z��q���u9���֫�u^$�W�%K�`Q��a��+�NQ78�w�	�� ���������J�M��/Z�ʨ�e��n�_�ˠ\�MQ�C�bo�ju��l��謸M��)�V|��q:`9��?��DP�W���~"�Yw��0!�DI�kͽ��s��_��(w��]�BŰ�+��,@:��k`�Ӯ�ڜa�˅�Ս�yOf����x�~�f�=a:P`�[���༰��<J,o���/�D�uٸ�_c������Y��d�b|a��|{���՛.�<(���>�0�,<!�3F�G���%�@�P6w�{�i�q�D�z"`c��Pz�t	;
��PG�2��@rM���	�:�DB�%ڸF���>��N׎1���LHD�)i�~K��W}�x��(Ɗ5�Y�@G��W�lʨ��'�/2I��(6؃4�� `��$�aʫ5�?U��R/���P���C:��5$��ؿh�w�3I� ��	�*��LI�	VH�}u&��@�>z�"m?�p��1��Ń7���,��>��+�w��v��%�Ư�����+���^#�fQ�1��\BB��.����y<=��T�E���UU:�v����$;��y��8��	���w���E<�f����#�'����c&��3/H(g�d,Ӟ�W�oǸ������^Nkݺb��;�l�Ȩ�kW��m���7MFSR��zT�$I�'�p�A��ճ^Tr�T���iO�I���]5Z>�Bک9ӅVPC�\~�/mBPGQ(n4�Asp�<N�}��l@0T����H�����X晖	�\���\뉐��J�G����J$�;C(q��� S���H�2�
��ei,w��߾�NP�D�	��{\	Y�!3�"/V�T�s<�-�>�x�Bj�9eEy�`k0��z�1�X����vD(/�����PU�`�E��-mtN���&���rT6;ڟ����
�:�=���t�M��%��K���,|8�;�� o`Ӓ�Q�C������JW�FCW�f�Eg���N�{=�� @�Q ��R��d9�.���r�W������4��m�o�0[Y
�4�7�":~y���"z�)pVa*��M�=�]С8NxN��u���)G�o �$+mFo����K��a�aRu�#ܣ��`K��$Ҩ?WXd��E�>m�������$g:����La͎��I̺V	����e��j���\`�C��e+�,w���#Ys;���쥬/���v���<�8�Ƃ�&���K�Q �;��+٣.�>pH`�`J�,hʟZ��i7⶟������"R9b[5��֕孥�@��i��J�c,�jD���]��7U�	�TQL�9~Nv]��|��q@�&ı��Y�b����!�/7i���;��?�d��]o-�M�����vRP��-�� ��|7"���N���`�U��C,�/I�zu5R��Bmu���يg�9)�G���6(��i2w�@޷� c�z�=U"�%��i,m{Jh#�~[���/�����&�5}כF� 9�AY�v��/�b��
�k\���38o�q�ՠ	M"��L:ZgY��	���l�៚����ag��;S��x:R�N��2$c%��!R���eBUv>��WV���?m%�KIg ���T2��}���m~�F�mk���|񀖇� *'\d6+����⿍0b�����<t�Ѧ��D�{.p�	d*7���ػ��@s�d!Ǫ����,��g�tK���V��u�
i�74�[q�L����_��]��&�!��)���\��K��,KĄ��X�biP:�k�C*���$$��B�2��rBz˥g���a���D ^�"�Jp�琉��)���ڷ�W�[W���"��,�^�{r�:(k%ϞP�������Fn��q��7T2��'ϑ 0I&3�h�7ˋp/����=�p � ��ڛ��7���17F~\چ��
 ��9�5�7-�K�Jն����+E��@���:��`S�2h'ݍ�0Ȭ�	ZY������.�ՠ��GrsVj ��a�(u���;s��k��&��"�2#Ă��=�\��Hl���Ἀ�Si?���/�Fb�3�H��L�mG�KC��)�ay*�{;��+��Iz�d^����`j� � i�)F��(O[���Z�'T�����.�2J/>ݤnv���O^�� �ϯ]��j�\�_�U^2���,�s�w���ǧ�T�����֜��fڎ�љ�V���y�@�} :S�?������JC�ے�ж��?����#�\�9�)Fސ����®�l'��!l8	p��l�DT��[6"<̍��v�H7ZY�� ^-�U���Pp^dp�Qw�[3��U[�iE��⸩�bۅ~̨6��)�����>Ŷk�t�/T�7S{�����51���aX�Q���o.l�K��^!`�~	�kIC��Ǽ@�<iV�V����S����!*�8���"����ǆ������>��66���o�4�;G�]w��Fڃ��D`̕)7�sW �W�C<��P�V�����Wl��Y,Ⱥ~]��:�E���H�����B�$3#��!uݚ �e+~HE�ei]{����f�8�w.b2�>�J����|�Bv�Ϡ�.� "/�8�s���6b�a�����_��د�$ъ~�	�� �e��}����X��zE+�C:�k�%�T����وY�yJ����jQ簐��z9ճ:�%ټ;���H�&#�����47�qv�֦(����N�i��'�J.�=4J���=t�͎����]�����@�E���ږ���Dyyp����!�~�˯.@bX�t@���֧l��M�� b=8a�Ge�4�����1�/%�kcPT�J��a��#
��܉�M�ǆD���}^�����e�a�	���1��)"��=��ىF9�gj�-��g�wr�h�M��X�����cyC%�C�gGa�P����.�Fca��� �!dn��z[
t.�
c+_�����>�D��������x8��1ɋ@:.�(|4�݀�c|���Q�Z�h2"����'@�4�п�G��U����X���7K����������u= �XC��;5�����Ta����TŇGF�͗o�>70|�@��O����Ƞ�a�����2�'�YMz2TМI������c�ʄi-���]�yY����x�w�*��M��$eX0�xȺ.�Hb�-�ү|_QE�¥�z�W�Y��Gg/���r|��D�R�<%ǣ��Z߯�&Э�I�0��/0��r�g��t�t�A��S���R�W�,_�"�#�D���o�4������mW�:�1ȼ�b�%ͤ�eD� �y��g��:���*��h\�^�^�ҍe���"�C�
܀�+w7;a%�K���?
�j�����r'�Ĭz���Ԏ��B­�茽�Xq�:�9����8fxҌ�^�p8A��zX�K���x��9Y�ND��E�s��C�K����oOF��V�SF�_bK��t�0��렱K|��[b��XE$'��WfD��y�CR\It��B�
x��-�0=`�Dg���V|�=r�hn�a���|�D"8���H�Yx�%�*�e�R��+"�1�bo�g��-+�!��w�θ��e�'�dt���h�p)_�s61��� }T݅?�e�Ck{U�����S��u��d���.��	=?2�G����nQ�cO����I�J�"�د�Y52I��oQPˑԈ��P#�ַ	��?���襬M�Ƴ��g�����!�/��t���l�>��x��dwͿQ������0+X�M���� �؋�v������u��9YA�S�$ty�����ߙ��"��b >�i�糖4�6��t=+�C,�3*�	{˸_<��ˍ��⎶� C/o�ݨJ���sIJ�|�6J���US#��*����@�����{�嵲�G�<��d���eiYmuoDF�b��9����"����%�Ö�Yݳ����4�$M�D�T�R����-�@�׼AT%����*����*����s^��Ɵ#H��R�Q��72�*_Cc�v�Z�>�3���.�v�I��y|�����g�%���&yL�����q�J��"�B#(G�����z��Y�)�hMM~��p���VǱ\��"� �؛�f�˟�g1�,1��3��H,�T�H��;p�;h^�|j�Em`@9��-��R"9��Lz.��e!�?j�*8��4���؍�HfH��G�վoվ��v:� C!d��݁k8�V�.��2b�r,�41���A%�F�}0v%���F+p��6�6F��ܳ��UfB��e��}��5n�=�%cXmzZ��*�N�imڮ�To�b.p厄���!quf&p0
�&�U�!�|�l1Ejlz�wS�$eA���δ��u���F���p��L	=��I�~0��\�]����M\�@�I�M�$�b�Ɵ۠�2F���#7ka�x	��Ss,���ǳ^f�6p�*��ʩ�9�M���a#���"���t�����,�?<xDsT��	ɰ�#40�@0���m���f.��Q�,|���x���DX����3�w��ՋVn }�<-7��ʽ��#RX��9t���r��E�Rݰ����x��+%�υ�d��=*�6ē����y���# vVH1C��ڙ���������|�L"���q�@��X
)�ѫ$�}aTH\j��h����r�V&l<��WK���-��&�*�`9��.i�fe����CY�����N����&5��SR��P�+�A6m�n��
$M}_�Hӆg�����Y��K�Ə3 ��~�J|��k��ۢ�@�����8�m$�dw�޺��]b�U�,�-��WB\)��n?��AUG>�w�9����1����x��6�*M	��e��j�?��і�f+��W�7�&a�#���� ��T�햅G�@{���xE�-����J�=lU\ee�N��6���rO�1]|?Ը��R\�R�[ƾ��UJ��f�K�y�����<�6ԛ3hߪ2*�������y�����O����S�ԈH_��@_d�����>3�)�2���q[�*�:��[{]�~'�[����X�V��\iN6#r�ԎֺҮ���e���gNV�?c�T�#ʭ��n�K6?#P�sÁ�!�w
7ӐH�Vaf��1QQSn �=>��ӹm�naK2��3Db���zn\���a6{9�
�>=ݿ��J1e���*{��|{e	�b�Ro�t�[&:�"�=dN����r$�YE����L7����#Q���<$	D@�h�&n^?�1އ+��!�t�T�>�qӫ�2Z�������(F� y�	po�D.��x1d9�.�Z^{��|&�돽�> Q4G��AG�qK��k4ߏsӴ�E]�i�^*(sщ��7	��ͫ�q�u�i	��U�6
+|����	������%n��@L��щ��1���|Є�d�J^瓿,�aʛ`�i8\�N�u�Kk��8SW���
ѵ����ؔ�'��T�~��h?&Gp����Q�6mI ���^��e������d	݅f�Q���y.m��V,=(�i5�}��֑6���v�S�;@��	�n�a�YO�=��>�˼��=*���w0�=cƩ��ަ�^��}�E&��b�r�`k����A17yR�Ai�;��v+Vv�ͯ\>�G1@�#K��
q9Q.�*
3^Jm�(*�3ʝ��P�X�Kh��O�p灰�tb M�W:�u�$��ԗ��Ӏ�$ċ�W?U���N���Ɩ����ݭX�� �%��>M��z:pAd��]�6b����3q`A�6{Q= ؇�y��j0�F�'9��>�&�lsf�pfÁ��C�{dG�� c*|��,��<����[�������&4�NA�^O��{b��(h4 �$�]9Ї�};�Pw��E�]�{�b�5�b��>tU����)�'U�H���QK yɚ3v|d��B�8��0?�,]�rc�����8�B�y�,�<�,��Qi/�rM���%k&�E�=�����㾯���g�\GL�s�@�=��c}u�p�؂�@"�Bfm��F�����oI�ڕ}j�Ǘ���f�@�ϛe��+�6FI�;e���Q�0�jx��|�:=�Ⱥ-y�Z��&��5��c(Z�x�រJ+�T��X���]�A�ƍ���Y�Ia��6�10�OO[A���	O0l�?ٯ)�
A���E~�;�Q#��P:�`�K�#A�(>�>��3��6�M:�3J{ʕK�I��d���(y�C;xB��w�6����.�A�>�O+U$0�s>���iA�l����>�:����S�!�#�y�?�%at@Q���6�&�������IwT�K��/���{x�WbQ��p��\~�b.ؖ]I@���M��Pr��SlL~U)�f!foKև�4�J��_�[�>Z_�V�I� �?�x���%�XY߮R��7��/[:h���UH�ݬ��g^�3۸5<X86�Jo`�*�m5�m�e�r��O�9�����a�Y�����r�#��2�~�\ʑ��.?��]x�%8D������P��N�˕�=���r�' ��C^�9�;>g¾�unK��CL���^U�
s�%[K�ef�kW���!��p z˯e�Ĝ��u,�{[C��3P�H.f�MQ�&���ȹt��	Qo>C�ϯ��3Np�������t>���!P�p���P��OX�;3X4���+�ˇ
�5������1�X{��e*B&�0x&f�{�h��lz�����O�W��Vl���>�:1�§<��<lޔl���Σ�3h0�L���J-!�g`����m��1��fv��a�<��9v;���<~�UK��kУ!@�=��U��";���I��v�ȴ�g.�φ�I2]Ey�A�QVy�U��⶜}7� ���17.D']�\6�d���Ⱦ ��?�_mka:������QE�<®	N��ҭ�G��`>)��j�u�� ���U���y��ŕN�k������+��u��k�]4��5��3�oO::z��$��� ˀ�F�~ͅ��d*�jd�d,�.�����
��L�^�
j���Q�)K��~�t����o��9o�n^a�D��=�L~�1����`����s�T�Z�I�ØK\�2ۭ@��H|Ջ���d;{{��Ü0��PE�6Kǝ�Jڝ�C���ce�� 4�E(d�3G�ZT���ro.\�X)4�m�p.�x�>tF`�)�抎�"���`w<h+��nĩ���[��+�O��2��������iD�8I�0�m��[�� �΁����,�B0i#����Hw�KiR�N&��7�O;����(r�P�K�$�G�݃�¡D��}m�o������ ���
������`�����q���K?�A��Iq\�1D���kf��)mr�s|A]�܅ob��ӎ(�ў��^"�_D�B\)��?�My���ПN����n��m��r�%"�X�,Af�A[�5�z��{��5��@3�`{�T��n��!�t(�o3ǒ������w���Q�!�B�����r�뤐(�|�oO��ź������i>@�x�c�S�;����͐ktk%��j "K�j�����w>9��he��*y�Q`����Tp�E'-�Q�8��w�+\J<Yuf��X�������J2X7�����;_���O	�91 �� �.t��9�y"���ۮ���z���|j�G[jnڅ�	'U��Wà`}RJ�ߘyOd��'br���~P�,3|յ6�p���!�DԦ�r�����%=u��:wCZO�P��FH�߈t^gK9����H�Q�����吽�b�b�it���;��&n�l{��U��{$���뮛{��"Q�joz,��3��ۍ��,��/��b�L�QO�P����=�FUC,�XĤ��ź1X}����%(���W��Oy`��r�l��1˯,whw�S��,H���=�'ͳ�
���ú��y�fS���簏D��D������}�t�o��1��-��};�),)vۻ�l�Z�ANX��M1!���D���8��f̧e�F9Q�k�-����b���nC�e������m@>nu���1,�4荋_�D�S	 |,�J��]���4�`�y������U�m.� ��w�Ŕ_�So �*���x=8�
&�5yי>�Q�����v���!�Ls�/�'W󼀒ɴE-E2�2iKT-j!	�
�����~��[9��5��e��8+���Pk_x-��}u���+k������e�Y�5�[��%S� 
ˏ#��v�S� ��UBr��c��^G�pt�-����c�q��������z�p"fx/��O�qgSȠL�`���$d���\�b��{�}:DV��R��L���CwWF�")d����{�rMX�wY:T��2?eBF��Q%Ӡn���Ib�|�o�~b��@'�dE%M,��Ou�}O��^h���h2�yQ��K����pxR��c��dp|�O}��A`9ۛ_��]��|)��1�)\���4�����o���Q~�1�,�Űx/ܜ�o�#�=�+k~~m^�$A�\	힪ԤG1��ݿ�ߪg�^[?L�nk��I��y��/�1�]p@��	
�m�Ne��eR�z���Μ��T��H��i�FYe���)O���Hwo$��$�s���/�iD&m�d�#_FO���v9�31�i����A5�������]/G������y�%�FU���|�e2��K{�>gn��>��=�N����eTk_��2PԨ�R�!�l����^��*m�6�2���Wd�1�N��7&��R�:�r���o�JоPBl+��y�o�������dG�E:��b���	���a�(�]4��bη��-H[Ø�K.V���<n���<��\5O����	�B��o`V��Ȣ��_*i >o2�=4���h�je�>��,����T�������*����@ɑ���J���cw�� �4���)4�p�]�C
�m�(	$`���;����k�/���Z&� �~��nJ��|�܅��םEH}1�{b��z�i��O����rݐ�J �q�:�HJq��i]��N9�tt��h8=Q��f=O�M�G���Q�w0S��[��#��;�u��Lf;�s�S#�(f��JsG�}���]F��{���Y`օʽ��u&��������	��ł�B���ߊ0_Cʲ7~9S�d?{��yK���	=����>?�� ��+=�>\
[^c)��MM���#���\��C��<�P���DP`�3�.J�S+���?��Q�X ��{:���U��f'#�O^���F��B�٨t��y�1���U�j��wk��}7����'O!]��j�i�l�2h� byol\�lz�Y$$��7�
�:��� ���:3?7�;�i�����
@i�ޘ�~����(m�D�V�u���-g"1Q�]�%!#�o͍�EG�qH��>olnس�]��LGc�hb���-\1T�G�h2�nW��`���V�[h%4-��׏`L�#X��y��ݗ'�@٤�.���t�k�������晴G��-���QL�=p: ��mκ�����*ƴ\.-��b��E]���9��4��.u�6�:�Ƨ��&��u���G=�~��v-H��{���=�A&JhN^ 7�|�]#�͸HӰ��<r��nV��X[8ny���A�0ϒ-��c ��SD0��Sݒt2o�Y>胻ܻ6�!�l�m̺n����n�<���	�(�-O��F���^�B��D7e���>��_im U-�ţ{���ob�^5�±��sǷ6�j�[�졌�,�~����h��I��ŮOI=o%�DbA%1����h0�>�+Ԑ~���=��mps��ѝ��j���Oy\�æ(
��`&����P�����|S*�C���N#�♪y|�k�*�!�F%�%��.t���(1Bw�h�۞'W�MND��%jvi̾��a�v�r)����H1&V�m:Կg���C6�Sr�2��F�z9bYj^����r@�,y@��Gk<L���IXa�P[�&�Q�}02i�2#)�'B*и��=�O@�R�$���a�ײ:<,2������2����� � G	%���+�w+4����r���{i�Ǵe�+!-�k�F�A]�0�ն�&v�; Do�2�^������*���#	p��+�&�?����H,z�W���=oU������Z@7�M3D��m���-	�&���}�つ=-�z�p�0\�\2N)Ck�fy2?�TK�綋��q��"Q�;5���9v�K(瓌߼����>ÍJXI���P[0�f*8"9��YCM��6IE��t���� \�h���B.�]������k�խ5��ft�UC*nI�	YD��-�Wrr|;.yv�#�&�?�P�w"H�6c��i��XR���_��:טv:��{�:1(�gF�jЖo���e�+��YG�N��Z�ؐ�si\!V#��Q�K{lO��0yK+����*�ܢd��1L	�mH\+��_�~&ٓ*y�N� �E�vp�4����Zs�}����v :-�=��a��Z�`��i�SP4���ƛ�C�<���s���,��h��G��!���or����0�;Z�&'���I�o�P�*2��0�G������C\�����J�+���b�
�����`J��X��S2�B^~��9z�U�@��{��O,@QŻ��c�Q8�6Ҫg���嫴
mXg��B,�,(҆�AH�kD񘱌ӫ��R������#��Ao�JMy�,O9_�N�n���o@���udW�Mn�O�9�8�E`�ߖaѥu�s|9�Z9�^�gK���ɵ|�ch�:��Q�A���e,�[�LiW��e?]*Ѯ����p���w���N+π�*[&�!��ڀ���Ȋ.��<��VL����}�>_]�Iu%F�sf��WN%��v��?�%4)��يƤ�J��*A���$��,a�s͐,DU!i�D9u�NP���.�����X��vPI!m��m���b��vP�^d
^�Ǵ����t�~}�����ܫ�<OM���s��'��`g��ߢb��I��{��~**M���G��I�2�N��T�P���rm��9?X��74{b�,��v�����w���1Y�%�۶{�h�SU�C��6"ի��:ۗ��؍��H߻p�ξF����*��V!XCmm�_�����ρ���05�6�.w>AMRS-+��.By��1�Y"�EZ�1�Ĺ����U������"і�b;Gοyr��r�Ɲ�~Ŕ �Z� w���<��h�]z�J@��\��zxIs��`N`;�o˹��r)��h�:ܬ`Q�5J|-p�.I���_�$� [K�{Z�r����y����b&�[
��[Ɩ��6Oq�����]H��>��J��4�k�s|�J�Xy� �d�����>����n�Y���D�3Y�f�QJ>?R/�:����!U����ɓ�}�U/B�T�e}3d�>˱X��Avq����[u�X�+�j�{m@=^��IZ�
����E0�����S�/Sd��,d 	5���^��������M�o,��=�a;8�s!�t���7M3�X�������y.�b��H�����L��~�A<�=r  �wW��)��]<��$��-�L�H�!2���%����$�+/u"������(�30��é��*l�J�����j.U�v��~��Ski6*���[�C7ݗ�Ȳ�
�����ؿ* <T��ֱּt�ĸR1����BY���;5w<{�6��Z�,(����O N���	����i�[��ݽ�۫�`�yd�t��O�\���@|ǉ_�2c�(���OKb ?)���hh�t��fe��Dl��]�����v�B�z�x-�������i���&�����D�����d[Oz��E�D�?ՃX�.�Z�b*y���ɮ��o��':t��9��VH��îO�c?q9�#`�i�o�ܾ�ns�<�UG%溛���#̕��R������Z�7�xnPFzWW�4ӿZ�8� �?����r�YeY��*]�F��#��쉽��c��+&8���E@u*��&3��+zj����Qf�_�*�/�pY�%@nv _�8C�{hi�S�8��y�0��gݣ��Qܱ�U ���&���g�1��PW��hyk�ke����� �ׅOk��B>g>(O��k�M����~̊Rl�N+��T�ᗓPJ��XQC���㻐�\b���.�u��X��"�*�i�vE��i~?����j�jlꕭ����d��\k��a�x�F 7.("R�s�^���aR(?�Ȫ��E;��lz�����j�h�{�XyZi��œ	e;y��$�7S5�^�B��b�G\�������)j��Ҝ���Q��]l̕ فc�g!���#��͉reX�̵�=oɕ߲��x�J��T���'/d��6��;���7�̶)���3�[c��`C�U�O�G���1)�G}S�3`�^U�f�TFNղ�l.��0N*�E(�t�f�iޮ��	�E��~[|����l��� �LM]ڤ�v��.�;X��׿��'a��7���CǇ��&�� 6RK� �� ���u��x߼�}��� ��ñ^'��C?��Yj��Jջ8NY�q�O'���(�)6"�����I�s.���������.�Z ~��Լ�Bͧ�՘��\�f_�2b�G��!���X��?,d�kt����Q�D%':΍uA9	D�/Ǩ+�G%J��̻���'˒��pE�� ��&����b�XO(i�����Mמ.��@o��-��@��JC�1�Z�f�*�����{LڒN��%�Mn���$��Z��m��ܝ:~'y0��K���2�ΔM�h�~�^��	1��ϳ�*�q�ˌ~=����^}���-���-�Kq��`*w���9ڳ+ۉ���A��u�2��ۭ��&ޙ��H^�ڤ0�V_yi^��V��`�����^Y��4P���J�a�ڮ���e�N�������;l5��Ѳ��إm�lg��EM���\.�A�#��ͻ.�s�|��^X1���c�&9�m�W��k�x���9i�j�ȓ�@��`���?�	w�ǛN,�"t��x!��Xq8z����.D�0�?b�"�1����sW��tT@����>����$ *�M�9��R��]�_?��l���6rj$r�+�� e���
א���+[*�`�v�7mL�GS�������cd��sq�?1�������z�Pٚ�y�����{�__2�(�r������v��Fz�3�i.�+%[�L�����жLb�7��2��ݔRݤ0~�;�zI���v���04�GІ�}�=�Y�>ڥ&��߭ʲ��<����SN����⢂�M�v�e`HͱpC=�<}�?���ژ��!�����|��yeÞ��`�`˃Gp�_&Z�KN���DI��v�Yd��(k��8��O���<�xXZ���	r�'�5���u�l��۬���@HS4'e��t��D~N�@�&�@B�U��~c���} ������{1�;�g��Đbqr�hc80�/E���uc���/��s��hᩑ�AxÊ08Gh�{�)�_4�>#E���nO!��\�3i�ܓD����\���>G��h '� ��R{�Nm���z�e��1P�*��Ɨ��MR������ݧ�>�NhU]q�a�Ѱ��?�V�/n���D5P%tR�HZ��/zn+3#5�/���͌ǉ�z��a���ܤ˚ 
s��aC��rT�z�:ʥ���E���J7�Q��>6�Ҧ��6���G��(����>w-ᥚ�|2$��L~���M���8�ԣA����.�P�~�L�J�7���q�0-7�g�iE�*!�~�M�#�Y�vs��&����-��0�$��u�z=��y�����;�~,���*��p��>���*���ˏ�8;�>���v�9�AN�$�s@,�ki�l�4r#��㤊�<�(K�W���5
M�]C+{{?�/�ןr�,b��^l�S{zd�B�q7wW���ռ�#���I��<qtv�Q�ʧK���h�Κ������M����n�%J�*�Q��ұ3l�`�g�� m�Xg��MZ������gѬز{9����x	��
��A`��i���|��c+�&�l�W7F����1�hT���]>h5(�I� �;+��\��?�V��cҏ��>�mn'�/�=@i�Ӷ���g�|ez>@˙��ER-��������� F�0�H�3߅�C@�ɫa_u��ʒ�3�
��=�A|�-�</t`��K�/�r'����$�[;���7���%l5ʝ[W�(�PQ�[���g9�,�]�sn�6�TBL;�
��u6ȹ����
혟��OB�G�S��4FһB�o�'>e�&������"������ӼU�!ыv�������L�8�Hio���C1r�&}�I� ��x��q�p�S��v�nT�$H�s�W��=0�?d̋_�9['\KBQ�"����ԢѰ3X��d7J�B�$��Y�j�2��o�T�$�;͝E��EEֿt���ժQ.���[�c�cy�����)�j/��*Y�:�@�g��p?�IІ[��~M��r��NoR�$PS�u��F�����,B����WCw�3T�K�o!!N��򿱪Z��(��u5y2=���� �5B��]:]���n��H�����foӼ�ۓ�Ē
����M��M�s�W���:����Y}7q@]����V!}Ao��j����!gOS�<=p[�w�3v,��2y�	"7;��k��Y�.C����� ��� K���,?:� -�}�8ߕ9)�?�Y�W���PѦ��%C���TN�Lz�5�� �E�K�N�KIՌbp�N�U�Bu�Kch�$"���̬c埼��1�Ǻ&�Y���]�l�_�'�ۅ�R7�P��Hy1��`�����]Q�պ��VUc(�xRWo��T�	l���tΡ��7l�yE'�/�cg��3�}}�a��o�i������B��lOY�%t�ē�Sɯ��
+]U��V~�Eu�
��X�z'	��'������Eh��S;��5F�4Y��\�B)��kѠ�sX>�*!��{C�^�]�NQ}��'��$˅Bln��/6G���V/A���T��~
E	ha#U�{~?O���|q�EsMq���l"�H$f1�ii.92)K����y� �]����1��H�ޏ�Q�2��%quҪT��'��X����������#:��hc;��<l47�SG�f�"�)����+�ށ��x��
R�	+�4�FP�R�d6�X�7�%L�2A�QJ~��w����o���&���
�]:�n���_�Bះ�Tj2���V��=�I�?�*{�_]̓ ��#Yt�_Ov��I�K�ì�A��X��,.T�߳`�o���jk\�Z@��I�CX�7C�q�Ch+�H�vK�_;;�L���&�D��ohn���a�S�"�A
$G7���f`����J��l�̂rJ�@���M�١�˾�s�GN�hRI��ex)xw��nQxA!>� R*�.��O�\���=�i%��Q�¸�I8��������I־�;!��K4��/��f*�UV��u����LD�T)��v�?��^����ڲ�F�Q�[�j�x�$���ma��=��(	/o���1�%5�7������N}/���_�|٪�俞��������h�6�×l�1�Y��>��D��;��+R�C��2	�GT�.����>2�p��^�|���$2�Z���!*��|�Y��=�5�)��5�W�ٓ�b�O���a��B��avI���ۥ0�����n��?^`�v!Z#"1}m����/<p�Ǵ��Μ.j����H1�ȯ�O߆b���]���p`�	cdt=���ep���Z|M�X_%a�e$�m]\!F�\�7���4��V�5�V�{�"a�~V��7ja��Py�ckuBh7��db�re�����3�L!�͖Q�W'�#��jy/��4�ӻol����Y;ܺ��3�n�����a[�6���v���2̳��.�F`�Yx�w@������9��Aq~�DH�:� �	��X��_Hh^B����"�&���L�ƻv��^ݿǘ�����1��
l��l�7O�l�9�r^%�����H��u�d���4{�	�,����Q�1�x���m<�R��/ ?v�u��"�4��f�}�S�⑁��Цc�x����񙚱o]�55[*Lz7�o64>+a��H+���i����~�4jqR,�e�?ΫUuLCн����W�M�t^Y�ƕx������<���Ho�Xie!	�#���K/
��������D�ncf�3�җ�Ѧ��k�$��_�_�ן�Tx�$��آ��>��ݞ��H����[��kP���\��Lޭ	Wb?�˾t*W���p8J������߳�K�U`����
Z�v�Nv�&��֤ӏ����Zpx`C6�`���~Fmq�T7�PX.= ��ݬe1�7F�_��&�ь���������E�։[�h{V���4�چYĨi�% ]"q���+"�K��Qw�Б]��9�7�1D@��[�2�M�}��aǲ��M�;6�?%{�3��JJ��*Z��jܕ����QK�
�iޢ-x��v��S����.�/�#�l�D���z;�X�=L����U�* ��pii���o�m�@b��y�����=�Y2������~���%tR#Md٤���dY�>�\�n����n�ϗ�/�9b	��w���U��q���̺���jB�T:��m�,!y�Me,ð��1��NO�>iA8���8
�-P͏޻x��D�p�9��-�3n!4����<�2���e�$�xs��1��
Qʳ�d��B-��B��{�+����T�t9�E��d�4�ުI"}�2�c-M��:4��VM��/L��6�M�_<z�1{#�ne�S7��4a�x?�a��h��{���Y������Yĝoe�C��EP��V��]?�D��4��⼩�=uV���;q�GB��W��Z:|���]��1��v��rp��$B�H����۝S.�+V����vۖ"v��2����:��aj�v��6Z�3E&����l��[-=�w����=h��UNèR����f�n���)7`�֖Op��S������V��JnI���&uz-�a[ͼy�˫ ��эYJ�yG�����fP��5���	z���Gy��IgT�:������՝�(�HIe;�]LK���-,�����΀'�m=��.�=2e�' �_K,!$+B`9�ɗ5���<�������Y�����Í�հs�$�+�]��s��W�}��0� ���nEn���E�q���_q�7iq�f� ^U�4�����y޴=m�ւU鳶��j�L���G�0�e�1�/c;�3H�C�^�tNw���֞f����5ܗ�,��N.?�)��>������ނ��xM8�4̔����U�?P�Y��%5�������6�վډ4�~�Y��v[e~5�3|��?5��4����j>��@�B �Q-u���3Œ�����s%�֐��P���5�� �740{���ؖ���}�v�,"Y�ۯ^�Α��W��1���l�4���N�UM����p�&�d���-��xpk>�E���Dܹ�,h&�G	6�5O�E
;�j�a}r%j�S�.;�ÓXcfr���
A���E=�� �U�{�1N��5=�?����2��TR`�/	��ȗ1�D;y�Ա<���-�VR��L�"��m��)��*<������}`�\y�x�� "i>a���U��I'4���2[;�C?�~�tvY�q�p�[u� u����)
*a��"ܐ�M�� k���	�-϶�h>�(ȫG>�� 0oR0�zU x��}sDK`����b�.r�l�f7Ž?H�B���?)�PNJ���K,|�9E��Q�ך�QuQ�\����T��~&��`�X ��>a��1x���i�����$��cB�t+ݝ�ߴC�D�ۭ*(�)��/��������������z|Q�Y�+���$'V�:%�hV�`�yDۉJo'ɼn:Y��h�a嗔5"���;6�a�������d��*JY�t��0�e29^>b<&���C��S��Ƽ+�+�h��)����۞�'����	�:Ot�鸳���C�Z5�*�F����D^���$�Ʈ���o���t��"I�����~���T���%�`�mչ��&dނ=����qp�V���<�|�X�'��ǔ�|מS��ʢG�+Bξc�4�8��n|x�s�p�'�������r�#�`2T�0��6 佈n����z�ۼ[߻ĵϵv�H�-'����k�[tN�o�峢�솣�?x@kN�c���/}�u)@QzA=	Aiԫ��~w� B*A��7��Vmb�t��\��#��R���jt��vb�����a�G���_	VԾJ+eF��ř~8���F)��>gs�������m;��FҸ���o6|�s�����׶ה�=fl� �j�$謒+�~Us��.��j����1�ipH��#=�1Hs c|�zj�ny�rMUa�<�˜i;�T����&p[*�4�=_Ǻ����grͲ�-q;t�=�td8���K��M��<P�f1+�"���pF�y^���x)�fR_I�r�	���N�V��C"�H��TRV�U�-'�l'�?��%w^�M3X
j�I��هP��@ϗ9���Ǉ$��Y��_���6�="=� +Mc%:�{�yo���������  �19t���[�y2p����o]����1z�rf�R�{b�I�ɻ�+�� }�E�_���2��J$N�F��<F�.*�u
����y���g k=�I>��Q��c��T$_�k�RM[[a�"��:�]=�*��B�/��,�*fH�����<�%E(����\A�
y�X'{�4�}�����3����$0��5@�CH4��OG��n&����i�^`n��>��DK��A?�i������U)M&8<��fZ��n@�_�?4�oO^�c&q�.�w땂r@��|��#?�6�7��R�A�y]��9�V��1��D�c��y�	?͚{�|�����U�A��YYr�u��:`9=u6�Y��'0����I-��p+A�C��󾩮\�d\�ٕ!�냛�v��(�,ǥ�"�������)��:y���|�uE�|F2c�ᶎ�eu��v�"x���|W�}Vj��NǸ���5���FR%֑�����$����k���aC,��;.����#�麐�H����ѳx��7X�9�Ԁ�e���4N�c�m�W�����5��S1�p�tl
�Z�GL'LF��ERz�-B�)�FO5&ڈk��j��&k���'�D�ܗu�&��ҽ\�x�@�䅑�p�*�q�!��B&��5���܎H!���^�랜����"�i}Z *Id����Ae7�{�#o���i����O#<����a�Q7G�Y�f��ksA�������.#����`f&�E�k���K��[Yw~�p�T������_�'���~��L*�}�X���W�Y�0\�>�n�+M�}��'����޻�jj��K=�;�)O:�Q�N1�Y����'O-$�ՠ��#�� b&�xՎyB~��]�0��G璶�0܉0�l�1��<�6=�H�	>Y�XX{>�Jz>�P�hP�>B�wڰ��z�?׆
&ҳA�Χ��+m˾B�J�a�28�JRm,�;�O��g�3������Z߼��e��z�����8�t��&�1����;��t��MDpۼ��Z�e����v޽��+�-�/�����b�S�Sؐ���2��U\��߼���pU��E{CrX1جD�|r+�/i�oþ4�$��2�k�lf�!}���R��i�u��-�%��E� 5p�H�ۭ��2��e^�W��,/�����GCGf|�����9��{M��'m�E��^nw
�nB�� CE���Kb�*n���_ܭ�Z�$F�ML�D �V�D�#���	�a��=�d�8�Fw�kH
�*�	!�W�y�+�]6�|,�n��\�ڨ'�!�'+>F���z3���U��EޢPk\��gaʘigoA��Ocl7��+#OF�Hy��"I��6 �h��1���w��5�J�$��}{w�L��K$݆��[��G�]OX�R��jVj�cyX���y����v�QѴ��
��
/ �4�B��A�Q4��׭��E�8�%J�ġ
w��x�Yt�N�i�F�{E@�?R݀:�A=v���ې"�F1��Q�����|JrR&�t�u�^��d��6d듢�|��g�Y�@��o����r�P��QH��Yt=��
9����n_�D�WЉ�����۬�N7!���-��Lj��%෵�l�n��~��n�F�˸�UFׂ/}�8��vwi{m���Y)����|��S����r{�i6��nm��D>���;�xyR&:�v'1$�@Sͷ�@�4p5�9ʣX�A�l����#�>��H���2�� �v6�6��S�,��Q�y������wm�z�ِ[�Yr*��D�����BWԔ�r��>�6L�Mp�x�Cs�����	TהxGO�(3�6��2"���Q��̅��D�Ɔf��^�h�%�u-
��t�m�^��U���u�V��X�`�}�r�5�������G�Fw�#+��f�|���!��@�B'*1ٜ�҄~E�5��D9���6��� x���?1Ya�nE!����p�&P1�~�j�!g�1���*��+GAn��fV��q���k5�$m��k�m����M�~I<������c���~÷�]k&T)�b������w���/��f|���[%��~�>��x�~�T��55��v��0��P���Ο&� ��x%��y��B�*�tW�x�p"fxdthT4UfƉn������al�dN�9��j�������Xa�V���r����(���X ���*hF�"�sfI;�";8�O�u-K�NT�*��Ú��m?5ޯ~'�Զ�� �
�!h �F�T�j��_��lG�,d��ξ��C�fœ2��"13��pP>�Tpozg�(qq�d����h<8�a
J4�����<Xw�NּRz�k:|���)_���-SE�{s�@���3"�h���&�"c��[����N����Л�����&�Nӫ��+I���u ��ju� xg�>A	0���2�;a�5�#���*���K|�*��R�ۃa6a�5��ɟ�D�̕�e���سtoB>a/��;m��������Ҕ,�l��OHuX]A� Ԟz��'4�l������C�XqqTŎ�4>�i�:��
����Par��cن)�w��ٯL8�j�WB�=T����X�`��6!`s$��[v"��$�4�GAB�H��c�=�m�Pp�A��G~��1�a�\N���_X��A�x��X��g��(�"���d�y���c���b���e�Y�?>��_bΘ�{k��1JFǌ���|��E���TW��S.��H��T�a3�{��Z?�e�E����m��(���6��"��{4��~>�"U�Y2���o9�N%���)ej�(�j�2øt�߰FM7�vj5���������p  ��=(��������pA��t{<�@��)Y��`�vz�,|�mr��'z��ᥔ�<W���m}�9��̹O٦����{%?y�.���&�JV �D��",G ���뇼��@Bɐ��`h"���=��t������݉�WK7�oӓ�z+�)��
���[���ȿ�!x���\�j)��Nd�n��ݓNGj��.<v-0�S�x���yn��\�&H����;Q��{F.p�Q险0�I���G��ר��U��$���s�n��g?�c�厧��Ww�X���l_�ȧ��<��;a���p�� %j����%����
c���52l�w���,��1ǂ�~�gIa���ӽ��-�rZ��n-���F=�2��!����-�3����g�B�F��=!�D��ɿ�5�."_1y�xۏƾ�d'72�d�7�Z�_���c.�i���qJ8��J��ba!�^�t(Cyc�tx=����%\�Glo�<ZTurrg���ʳ9�ĭy��
<z��r��<�����s��NN�x}ƿ���ʶ���'FE�-�����:�@�/�?ӧ�
}!g^�AHu'����+��f�z��!+�z�N>C�H�W����6� y���/��[Uv�+��#�6\}�݀�G��}ڸ�59�8��4N� :B+%y#G��Sm�?�������tNN:�2���a�v�n*�7c���6���&'X+Z;�te;���r�Dq�(7�,�*r����~bv�*s��w[opP��<�`���	[��U�����y�t'%K��v��*�����a8L^���
%�҇#I�z�Ӛ°�6�����g��4�B�i��C���]�G*��R%�Ox��RS3�X���m�e*0�@I
N�z�d�R��/���	�;���1�O��1��a(m0�d��9��^ƥ�̋Qqt[����2GR��e� _�f6����,�#ۓ�4bx1��E+A,l�Ĥ͑��o΀��$>gO�Z�ͳ�5RQ�,;k����A!@ӱ0���wC�s^��¹ޥ��+w�`T����5���Ȯ���B��#7%� &���ɦf�ȣj߬�<2en���r��b���{:V$���dv��2X+��/N�Bj�:d�ڃʓ�[�m�~+$���R����-��W�x�))G��Z�u���y���U7j8��<��*/��:.ؙl�d�5���ȥ }�-�٩�R�:���p\c'A�C{p(��)�9:vj�ɭͥZY�W
Θk6���
�՟P�_ %����`�����7)ͫk�T��¶��I�ǧJ7�Z����P@*�wJ�C�Bj�"�S8(��]��� 0%�Ԯw'�->����`AaT L�����	���e(�`Z�ۜ�%�0���3;bҟ(nxV{��]U���D��5d�2N��ϼ+k�&�<Ҕ�M�@z�O�@1&'�߬?���	lupwڢS�`����!z�$�9㌆�<������P�� ��3�8@�4}�{W�%��F��
�<�t�Tq^���x�El�9��MP�^��m��)N��8���
�뚐����5i����dNVe�;��u�mA��p�kBD	��C���H�g�U�ۭ[���PU M|!��� ����rQ�2(3x��l
e4;8��0��F�_-H�Y��q����R*�I�36J���6�Dn}ʦ7��~f*���:)��T�ɵ3D'
�f�3a��8��n_���L��`��n&�,�g>Uu�? ��U%�\���s=�v�ůW(s��Z#Bb��������>q�o�B����'�AP��t����[.��� �f�^B�I�٩��fLnX�����<ٽ��v�I��H��R�vU�3���~�J�_p�����@�.au�s}p\��@��ʖz���{Q��#��ش#�l��ϟ���'3��姱���,��`��A�2��`�o`���bC�@n,'q��M ��,'3n)?슝�?l����]�Ѹ ���O�'����:��=�k��/�|���{��7���:��|X�t��8?��n#���P��\�F*�ܡ��A��A�Nx���"��"ȸӚ�N�.#��׶�0�aMT�����WwjB�rw�w�$T���f2���3����+������NX�K�T�tsҖן�.#n��W�Ņ�5׻E�	�15��G�bw��x�E��Z�U�PpC�[iAݘA��"�.{�y�@���5�7����|�v^$x���2eE8�r��x�w4��~Șqݱ��max;~�	h�m�Q�U���Ć��ހ�]Jҿ�1Sf�ll`(, ��**��I4�U�tgӭ��+�&5�'��.up�X�;�ԥ�ٮ�v<��g�޲#Od"S�u��ktU���X#>2�,8��@���,�ow#-(�+�I7F����y�I��͒��zn���y\�a瘆�� �ZV��п�������_P#	=����?tDJy���H+d��,ˤ5�"�š/)�l�q�
��ƹE������ı	��(�W�,�'F��چ��N#2!�#o��2n3|����`��%��։y�6�;�4��i�MH�`#D���Hg��q�u�$�K ���]�0Vݪ���3s5Z��^A����G��Ȣx�d&b��6�`��H�Y�3 �nf�'b�u�H`�� ��q�t���:6�������f��z�k}���Y�SΩӗ�T��'V*�'A[�O��wH�KW��g��5S'Gk�Kɫ��y�pf����7WB�������'�-�N���Dc��a=D�T�>��f�WF�!�ټ�\��4��~��_ъ�o����Ig5�^2|��H5���yS���R���yf�B��m����7�7�$�{�����?X��nJ�fz7:�Dy�2��ι�Ӡņ�k��Y�z��� o�2c$>���Z��|��I��L�BhB���kB»��)���>n�h��q�z�ف�6d�"���h�����3Q7J��7h}kDF�Ŗ��n�����薮ȕk�����n�GKf*�cC\E�d����j7{a��%�#������~�
֢��F�����^��Ψ&I6����^�&��a����f|*j�K��J������Lg���V�U�n��S��y�i4d�~r�8���D��ѫ�E��ǫ���'���~/5�5�����ᔈ)o�k$�F��ösx��r!HPYfY%�REc�vc4��:�G� ��[z���叹Q6X���=E��Gk*��>_�^c�`N���qHћR��~��$5���g[g��;�TRʪ���
��"�P�|�j����pp�&4���5.�L8��p��j}u�:�yB����b��F�j�<��b�,?΂})E%��|x�2_�2}$�w�� Vz��Qÿ�c�/����Q�+���D3t0��`yD�XfTA��ok`��e�H�#��g��&�F��+��7*�ř�h�n1=�\����A�1%�v-Y���Z�H�'�D9�EH|����!џh0.��َ̡���t��v|�l����-�\*���w�����"'���o\jF��Z�x[A�P/rM�8|�z$�:K��r"�����]oj���U��ޕXFhR[�"�Z�-���<��ᚙ�,�t¦���a�M���FO��2��Ő��82��νT�6�ַ������W�2�w�e����8J��Q������ñ�ՐS[bE ���<Ȇ�
8f<�n��L<�؁�s+#���9���	xEI �}���d�ӎb=mL�=���V��J��<�і�`�Qibi�3hZ*w�f���9��	����rWc�����ˋ����_��*����7B1�}���Q�)�2v����(WLT�=�|F��>���kD׵b/R\� ��D�G��"�l$�؛3�Z{�Y)p{��Q2u�䱬�"(v�4�\<
Ǐ|8�R��"S���Ms���X�2-d�t�&e���ej�Cj?�.9de㑱�-?�I��j���[em�~B����7���;VA5(8�K)<Ү<��a�[��.���ë;'��(�ps�*�s���\.�$��@�:~�\|*�8��^u���u'F�.�,�
m�pM����_��;��8д�/p#Z�FY��p<��ؒ��c�-��R�5��>����&Ɣ<�EVBE���fT�ٻ�;�
<ӱW�P�A(Ш$Q.n��o�-�oqB�v�f�Hԙƶ� �L��<"�h��2�2[)�����h�Pe*�a�M�?�,�f Ƒ���d��̬J�L�8b�x/e%��ޅ���%}��Xmi�ʠ
�;�6%��ĺ}h�/�܊.���Ă�oA�J�������r`���u���[�n�����i�;�5z2i:���`xAٞ!�GM�YD�0�'�Hb.~�M�[��e�n�
�=kn���yO�P6�E���u�gj-�t�+Rn�񭻥i	.��>���/ᦊ�<r{NT?����UV�����Ϊ��-	 ��؁.��_�����k�n����<﷬�DC͞�b�7+6����3UI��s��$5���������7�G\��z+P����k�?Y��z2r���ka���֎x~���+�o1Gq�t�=?��y��fαݛO `M�-�^���J6pz��]�GRN�Q[�'i�
��E�d�9��.��XZ�渝vh8ԈD2B�JΧ� ���|B�'`w��l�vA&�"�AXs��vWZ(�X�7_,1�̎H�uwj#2�m<��?SKk�Ψzjߨ=OB����w�k���P�2�1����L/E 寰�8Mn�C��Pj��b(7�q�ǚ��H��,��+�HЉGڃHFQی��>3D?h��]�����KW�~�'��Z�>!����+����$V4����4a����A��V��V���k�0U��߅ٱ8����F)~R8��:��f�aL^b�)%�eX1��K��S�c;$m��2�`�æD���͚�h�u����8z����.�����T0˱<�1��6�s2�y���hO���kۥc�-��E���~շ���0���S�Cƹ�}�HLq�%aF1#���}p���dw��+:���a�߿CI{�����6v%I�]C"�zKݭT蓠I���D�w��9��Logг����NW;6.hc̻'��?�s��������n/�PC��e���̽��w"Q'���`[�)�d���1ͷQ�ժ�D|/�٥�+k��؝�LX?�WFi�� [�@��؁^�(")jiDCV��Tu�(Y紳)䘄YJgrt?$� �t��Ύ���kB�G����Ţ����-AY�;dk�����q�檙�uH锐TX���ӻb����ZVzjf~	88��+�4Y���ܒ�D�
��u�����:����i�Q�Q�;tf��W��G
n�N+9�2�o���݃�i�y���sj\Z~���P�&qi4��^�y���;��L��/,Xad����"Ɵ�����]��õ;+�'��
�{U�`��b�ɗ%Ǚ�b�%����Q �V�V�� ;	�����s<���5�*8��b�~��k��w�z�M`�f��(7���߬n[���?��NDb��5���f�k1�[h�|@�=\5�@�6�!��(>��5��D"qt�$B���6��NM[�7%>���g|�V��7)a�������0"����#�l�A��1Ml�E�x�:Q�?n����G��h��3�nbۧ���_u���GP���M<��3����.<�+!�빊j�����z3�$�a1���W�D4��ίÐV˖��!f�����6uC>��eO:�$�?Ғ��*¶�8��8�+��:�6V?,��� �ޥo�(��rvq�5 ��P{[���$;���]���z>���H��n�-��6�����g;s��|׬1wd&W7��E��6Vx��:a�q11!S�q�G-~�/���P1_$�*u&u{��2Ue&�ba�YO>}Sn�zG�k��O��u9%N��֪k��u����n���1
vZ�M$�ɋ��6�����I�UkAƾ.��9(����QZ�o�P�J��N5LE�#a8x�N�kՔ>jn�:���������O����ʔ5'-[; �˿���y�F�G$���p����$	b�<����� �O�-C��g��]��>>�1�Sg��U"�utљ������e=��\�$�v��q�%�Zi<���SV���o�Gc:k1�F��*���Ƃ��R��谶�]{�ϏX�d�ކ�iw^�ϫ=�\l'}�>�8v �[���HM9�"���>�HJ�p�W���y�)����vi��?�L��vG�BP�H���h�wV��x��04��4s�����@g1��_ν�5̡��*�@mt�?kO�6M@�����3�N����<�P�mB��.{am��H�R�T��	���_��*��~'0v�YNat���pfŠ�f��v�V_0���V����EY�V�z{���Y$�/���k5w|��n�%�N~wj`���2��B��K?��t)$�ـ�:�N�]y��}�(C��y7�co���+�����L���V*��|�`r� ����N��r|��f䙩�	E@�jI*3b�`�g,��>��=6��6�m1�j)�t.P�)�?�<�l��6���_ρ51e�Wk���.�͂E�rZ�$hg����s�k��@��؄|:c6��߃>�;k�8�PV`�*,�RlE�[گ�����)����|/�\��o\s��,��M�O�����+�����+M�2��1��sp� ��x�j��S�u��V��yB��8�)�>�M~�n�v�|k�sVi�g����� ��D��׼�Kb�Ԃ\C l��f��~�����l�������9n�h�tR��A�ݠ�¨R��=�b?�C�6b��A�>�N��lP�t�G� ��+�����r��!�hq�Ym=ƨx�2	?o�(��#
�(�2q;��It^�ȅhQ�幧� �V,7_�pl|f�*{�x�z��%����yrb��2Ɍ��ǋ$ ���ZN2�I���ur,�����N,���[����j�� �}IǺ�ƣ9K���o�sF��i���J��Ou#��c|�ϐ�;=�:�4����L��#�^[[gO�b-��X0o!�P�(��]���y�� 1�lW�IcŦC�Ώt�1�ݣȐ�x�����>"B��j��uXG�_�^�)aS?pX weg����t� ̲��'2ѣ78�AT��B-%5˶T5��z�ǢD!c\tח��%@����^�5G"�yR>4L�.P�&����Vi*���v�����mW-nw?��.d�i����BQI#���]���s�ظ���U�g����B}C�˨���
�=�C���R
�M+��̼���wR���p�����o�	B!q�*6*���XtnM��d�Ů�I�]M�0�f�	�9�)c�*A�au{x�0���{�)=�s����h�d��ݹ����e?��ɐ�D��M�u��ʲN�XҺ��G�e�&�h���4����?g^ �Bv/]Xx �fnx�5�,�4�Qߋ�!���hUJ)�j6s�17�S���mzϩV[����I�a8^(ræ\��Gh���S: ��p.�@�^���M�bp�vY�7����O D3���D���;�Ga�_����|�5��g#@��"�7ӛN���`�ڇ�n�	�k���'�S� F�t� �	�=er(2S��%�����K,�Gb"1�zua���}��><�������*���|����)��s��fi��OSq=�����5]��u����9#�j��β���~e��-'j��^���/Z�Ȓ<�m����|����Dt����X2|Q4\�'d�n���,��t���4�5@�^d��(�U}�3���~�7I�q��D���qǃ��`���2�$����ivİN�v�q_� ��ޢ`2��A�GT�bW����Y�a3@���0��Y�h��Zr����k>�GLm�������{�;���(��A[�7�f�b�����R�UxaSM�"H��+,q��FK,�&]��\aa|��8&�J߂e$�!\Nmo�V�T���g��s�i\��2�X��MJ��:��cV>?��x��pk��2#zH�1"���V9l�6�@'X�*�@�k��:F�+1�0M�@ixgG��<q�����w��Q��d\a�?л��}�V�i�*��_'��X�,>�	%|�8�<�k�M�~a?�1�j��:�p8�t���6��#�h�J6�<����������g)f�Cs���L阶�����6�+���/�Ն8=�`�7=N����.C9N[����O�ػ:� ���tX{�p5X��Z�0#~��GZ'1<W�!Z��V���B��!�F�[6�p0W!W���$}�<�8������_���d.ef�Q"�Z�(<"�U*�%?4���,$X�D?]V\��1��t���l.!6��^���_�P��!��b���H+���n @j�ӭ?�w{�\�V��4N"�b��|CÚX�/j�ε�h�s��*�W`ȔO�=�B"_,�f����brc0|'��vZ�D��=�8�Bu��U#c�O�&?���ڹWj���J�����@�57˦���������jI��P��]Ò;�ن7A;Nww��Z�M?��梔����3FH�?��Q��UZ��2�I�16v:xK� Qdrq��~����`ns5��#�@�5��O���*;&]L�l���~��H�O.������mK�+��{0(;`�g��:�p�C:"�N��bH��\�Jf�C��((�_�� D����s0e)�'xK7i;���'2;�fi֯��4״2RQ�1��X/Y���-���V)�-�S1��Q��v��	� 4%�4��`$����OVZ��$���,����P������/
���x�@!��mZsop£��]LRb��8�niY��Y��
x��d�w(�Љ��f象�}:��GD�?�o��h�ڞ2�BƘ!��"% g�Bj,X!��+�L�D����%n�]�ZE��|7ߏ䬣�ܷ���N9>� :�"�o����װ'A#�Ĕ�Mb���>�(�N����n ��7JRs�~��{K#�IV�,�4P�a��������F���3�nP`6�oJf>��;����4�6!x��[5y�B����	���hE��͠I�`���q��t'!<Ց*JeQ�K�ʩ9��\X��1��-G�%+D�yc���.]9���b�`�} ��<�ǜR+�f�_�S���-G�S sW�n�	��F)�Fr_~ƛ"u�\Uv��w��XS��>��	 �m���A|,��þ��� �O�T�)���?9�
���� ^? Hb�h�~��8]�6 ���VQt~�fJ�ه%��M��cf\�t%n�İ�Z�zà�pun7�܅�h��3+
��&W��d�ۦ�[13�;��79bQ�G��]\��[�����L��b"��u���U,�(�OYq��3�\ӡ|���g��#��a�Q[><%���X���^�+�>�bA|cf�w�,I�! c��o��|�p��~�x���\;�Ngj9���c���f��Fϥ\���	�&�q�3We/����C�!���a1�"bI�G��;�w�&�Bo;D,��x�p�x?f�)��{".��ұuO���%.����/��fLg�vöF�,�
O�zfǜ�*���)b��ɬ_IWxACu��<�w)el��j������!]��wz��������4_�x,����-u[/o����W�����Y�Y�k)��O�}l�����PGi�}�~�]¡�aK� $�LBR��R��[��O�)�:�}��3��
��C�?����hu����Ԇ(�!�e���P'����u����&�|�Gq+z,���NV�2�MKuTc�[�Q��r� �$�
��@��1�ǁ;��3D�;�t�:������d����α�*�"~ĵg�[7��8�ߵv�8ءh��[#C/ۖ�ޔ'iq�K�|6.($���]^�3l`�N��Ψ��H00ǆ�")7��J��g��:�݀�C>>�5qC\Z�/I�<� ���ZT�
H�b�V�'}a��΋a�4������k�D A��׸�����Cb���x�I�����Ҙ��N�('h_����_�G
�K�����/pU��qAo#�6��ۦmڸ��t�fng�q"�'��.9�E������|X4�3���RA;G�j��^��`w��9n�7F���%	"GS�{�f4��˒��Ml��
)0sv"D%��S��EA�킩^�I�'��;Wۄ��u
��n�=����nGG�1��b�
��G�e+�$S��:#e�g�h>�L��1
ȵ�A�c�R)ِ�]�,,�DW�O���T�`#һK=޽�m� ������0�O�:��o�&��L��>�#�9�<�n�Tim�V�E�a��L�A�[������!��������l�������.���fϟ�3Tc+�E����#�,7�D]?պ�I�V���C3�t�4ו��H7�d��O�{C�c2\��/l�aـ헤��m铧�>�w��b�Bl��Օ�tY�,X��z��b�4�2%�X�n.�#̽"��I�'���)]��VV��Z����]@K���҈�!g�C�6��Ҽ{c�X��@�|n�쏕7`O�We��ׁ�"���$F��g��]�2h"�4"����G��=B'��ޞ��feԹ����zu~�'���lCN`S��P�466�Gi�w`1�/�'F����ΎY�)c��7���6��1�}�Z�kS����� 4b��L݄G��E�0ؒ� cԢ�Q�'����cI��̨��ÝMU����ݨD�:</�X��Jy��*�������3����R���w����  F�*ʟ5RsE�3�����Z�y��aMV��u~l0f5߃A{�ژU�m}�3�R>�"~C�,%������<]���7K�W�lv����O��&I���Ly@ǽه�d�\��1�lU��u� *��ٛ�A���*��s55�� lN�,���_��
���L��X��7B�.-�����׮�s��ͺ��m]��ԟ"S�����l滄V���w���in��p�.�74:�G����dU������M�����B�~�J��j2���ā�C�*�A9��2uU���^��$�t!X/)�,�'w�����'=���9=7e��uF�+��G������Wh��Æ�I���C� 䭛h�4/%��^�r��J�Qd�j���[���=a��|��w<)�Θ3=j���)8���6��s��9�t��`4|��9�a��*fW�����.% �%V��Ր�=�Swn�u{���LM�Y=�%6|o�1�K���8rd&:�i ADʣ�'G�c"�k�r���X��dl�O����`x���n7�pa^�un�qf�;�y�bcT�q�#2՜��z�ߒ����q��Po�v���ʀg�3�!"�����rT��Bj�c���j|`�����FBB�+/��3#Q�(����mn�)`�ʾ�T	�nλT=L�(կi|�2;M�;�&��~=������|����Շdv{�ֽ�f|��ՙ��\���L���m���(]L5hH�ܲHNi|�0�abB=�՜����A�!ٰl�UlD"�o�f-%��fz��6�,�&v����/B3���8 4X>�t�K8�@\F`ݭUY��]J\�� `-|������{g��*��������n%�\�\��y��9���9rA�Ԡ	K-�=�\�=�/S"^�nv����=�K����?=��3Ө5_�Q҄�۰�n�iO%!���w���IM�#;��悯�T��O�ux�7�z=�S�������+��t�=�6��n�j�,Va*&^Sm��]�T\ۈ&n��~3p��ڵ��Ag=�A?=��ȮV9<�]��b3(p)XgB���TfR����^H�n�\?-�E)OKtx�L�{��JS�$\g�P]ؗ�zmۜ�?�f�ɳ�-�T�;;�bp��B�O ��a�|i��,������A��T�Yh��RA�
4��l`��R,Ȧn����w�B�n��]v��o��uc|���F溛 ���2�j�"�>���E�)ݱ�GԈCGz�@ AOz� ��}���]�"���&���ME3%��pk6L�\|.]��X��!�p��Ɓ9�V�WX�{�D��T�)ޢ,��
4�<Ѿ	$�`y�3%A�p2z������c���9���&��/�M��� ��Ռ�z�6�x��3��tv�����8�P������ �9}��}־��2%�F�h1m���~�<�������<;�_������2�x�@ʘo�L�l�[��x2R�c�����m~���>�>R< 3�{�7X�Z�{[͈-�����-!�_,����O*<3���"D� z�Ԡ i�ర�zS9+� ���Crg8���
N+�DmW��D���������|���z$7�\OV�_�\��7�|4�ϕ疃&%E��A~�O�U��2�G 8���a�*np����NV���%�����j����d��q}�5��6�F��u�r�1���:Mry���6��F����	ZHw�)�	����������ӦC�U<�eȧل�����q��ׅ�:�*��g�W��>��P�%�Y�M��\K5M+���}�R^�`��3��I����f��1ަ������g̔,|��Oq��} o�=���e54���}���rڬ-� �Juvp���E?���i�� � ��"q�Ri\�L�:F��y�z�
��P�HLU8ƉW�\TFw�t��4�\V�|�;ϾDi:���28��q���?ĚUnE���+���\���}�hy�L�j�c�.�ȿ�ާ�|�F+y2���y [Be����h`�3�� �7��j[6G퐶�?0z=�ąJZ�0
˹�5:�*oq�N���>�t@�9�
c���ߡzL���U���y}�  `2� ��z�Ec:�JY��M��y��K�~b^���5�s���V#�Nq�2]�y����泿RS����8I;+�����.�Or�Y5�P$��eR��{`�t�����t�[�g��S�C����qN���Aޫx]�
B@�޴��y�*�s1y���+���l8�QH�E�S����8����P/n|�|+�;�%���M��
e?)�ǂ�hhMdHk��2�p�0+0�c��J��� l�Az;Bav�K��I^�_ЙY}k&d,i��X�;N�u�507*��]!K"R��D)?�w@4@t69�`�[�ޖ�s�cnN���z^ۢp�ҹ��ݩ��o+j�ʱYa�Cƭq���j��*�*M��	L-��.mD^HT�*H���d2�P[�{}�%$�Zۼ3�yL��ǻĸ����
����cNګO���Ѭ�!\Ut7H5��j���P��\�j�k]�*�dm��1����iE�H�§Nǖ���[�B7�����f�4��-"�E�1N,}c�k�?��e,��x"L���Vo@F���{�u%Hs,�s���uW�_g��*9"�0[�ق�p)2��z��f�,������F�J�ˎ�;�k~%��>�k,���b�������:Uj%��$*�j5�j�-��#�H��3���ˡ��,��f����ȍ�-x���i���S�l��߆T:�^	�^�vP���m��}���^<0,u0@���ް�8��'͆*î�`Y�(���:X��=p�2���B�om���o�%�S��	)Lq�"g,�M����6��lXf�-�$�|)��A����*�*/f�ɷ�l�^f<��eĴ�P���jǅ#|2^0.�����X�Jq���*��C�@���N���Я %d�T�~S�����M�{l�Nkۋ���4i��S������
\�@6*���*YT"6�R�7��?*ғϛf�8��w�XO�1=������g��9�W�K,s8I�m�cf8�Q�D���7��Nc"CC��nXY�����Y�����pd�p��E�;��J�hAE�3N4z����|h6�:ǽ�[�B�X����°�:�T�����Dh$���%J�z�e�	A`c
��*��{UIM4�ˆ9f<Z4�-�DGތ����~{d<cߝvDA�n��e����N�>=w��z�=�g�δ�8��Ʃ�7N�` �ϝ0f�`�����N��5G��ۊ���p��d������B�O�j�ޮ�ݴJ�H��|�)���cX��+U��i �|�w���m�q־d7<�����6c���)b��n���?�� d��s�����۾NBlz0�ȇ�VmɩL�	�Z��j0��R��%�X�~���gp��6�-۪�?���T߻&�����A���� �5�p�[~�"������ �C�m�p[c��84a�^b��(wE�&�{<�����u�k
�1n M��ᮢ>���0@"E��
C�:4�) �sFyp����m�$zR{}�=(S��c�*��S��
5ѥ���L���ұ�
PeGtu^�\O��6�*����7�/�I͇��XF�&��kg������k���ɤF������1�y|Jp���{L��Tj"���t�.��VkX�9%+��q'�v��Ke��Өȁ��ji �7��L�����d�u�а�f�w����B�Ŋ���d�{v�3�Y�
!�&p9�:9�{Px� ^Y�C#J:o�bg�l����C�7f�P��!�Xo�B�?p�T����e)u���'�K�Py:��dU��7�&'P;��j�FX���={��:����PL�T5>ԙu�#kw��x�=DG���&6�iTa�r�c%�+>�nD��TE�Ϭ��8r�����O ��~Yt(��@P�S4��;��Ug�l*7�輝:��%��+��g�K��c�U��N���a.����{Q�A �c�<p��́ޗ���χ����ז�A�Y�9R����/K�Y�N{+�u�Xq\�R(�~b�͠�Ѡo�I��I���TC�����&ʘ����1����Q&9<�f//�F ȋ$^r�V*SŨT����i���m�-r�l1��=�j�Ӊ���`��x;-�!����JlbjpcL�ޔ=����FGCE��\���g�PRK�}ct�ّ����Q �4�f,l�@wͽ`N�E�D�_<t��֙�շ��� ��d|�ݏ9\S+®���P���݌���w��Z���E@����䷔�E�	a3��[����#>���i����������`3b|Z��'I[�li�㶇A�N���O���GW�t;	�g:�sN���JX�#G�IZ�gu��i�G��`���!��T{�=��_!�L��_gϊ�6��Tfry5bq	D��cQ����Оn ����i�#�JG��<�B猂�P���+��E�3&��lo.e���<����K(���?�{K��0�8�bk�_'T���O�p�4"��:�-'���W�T�ɸYN��z^r�k#yt�f��7�]pJ�\����p��sX5jJ.
�ifW7��"5�i�˘ȗ�hi�[���ce7�n.�8%��=��"�"�Ov�)���9�F*A�m�c��J���%�����k����A�Ov���ه4C��� {�rqE,�F��+yqy��x^]�I/�(�3�a��s�U�/������!=5����o���g>nZ�y��h�3��Z8������������{K�Y�_�8;��Y�#�����vk,si���R���Az i������\������#�O�~*��Ї���x�ѽC��p�^[<�S�	�FЪ��/}�S�d��jn�&�
�+BA�[^�p�
_�,�����=b�q�
�[C�YXߪ���֣�X�Y^p ��+�;ɦ�x$��^�)q`+��:���oV�V�b"7��`�7Α#k5����{1��	��T��
w!�Ks�D��gz֝� Pö}/�[0Q�Ut��D�xlf>ʷ��G��c`��wzz�n`�ٞ�fXX�ؐ�^�X�Z�,f8����Hq�'�/�%C��8d��j$� z8ॳc�TQ�`��?�7�a�N�������1��8.f�%�ƴ��G���F~��W{#|�?М�b�����f٠,_Wr�,?�D�I�-L�8�I�7=K�櫑����
�[ �g�?���@��[wҺ��m�C�ʏΝ����D'�������[d�q��hy&��tD@4�x�r��)C7�e��RN�W�}D�ǖ�0�k��<v��!��g&���Y��4��ufݽ��~3/έ��[p�Ǹܲڲ��~�΋Q٣��A_�5��D��0��@B��d��^���s��̑K�<B|[�0`�#p�r/�U3䬞|�vKz6j��x��B\�	+/_�${
ۜn*����jp�+�B�pھ��J���mӘ�T�Wʈ0��J�J�`s[H	�ƫ��X��1�oq߃.�B�п�w�p�i�Ǥ��:{ذڿ�����SsZ����_LKj��/��}�H�h/F�]�\�?�2�쌉��f����s|@�f��d�?����-J�%*��u��݃0�(jɨ������r�{.(\/�#tJ���YB'�THt��u5�\�a>����j�� �k��k�d��W��������5qB�s�Ճ��ʰ�-+ʂ����ʡ֡´̈��I�y(��:&���h4+���V�ɱ�=#���R�����:x'�$��9[v�/�TN�?,��z���KW��E;2Su�-&{�<�^ҙ�":�DY\5w�k������Eu�wz���nB� a��>{�r��UBҖ|@�}�(EAD4��p�BRu��o�%2I�Mթ��.�e]�l�y��ܺ�9�}vp� tN��Hg1)�5�E����A��zl$�/��
�xS���.�%"��nyiUi�F��^�"��RU�����H~���Dۚ��ZQ�2v�Fa�]�zLڋ)��Am���D5�mzIʻ�����/�>��\��?E*֮\��E�m�h贆$�w��4�iU�Lt�~�l�W/���&��ƀ�Ů
��KRl7^Ф%�xg������u<�>x�K,[@l2}9�-��F�O���l	���DX*���ܫ+��A�#jݫ��;
��?�!ҙ��8wz�(�W3 S�����~^��T/�B�˻���=�񷫍�or"���FJ=�d�f%i	�e���j���C�:|�|j^$�k�DO���F�q�DK���%�C����T~���)Q�]mg����x� x�RB��s-:����
swc*Ӌ�}���N�l,�C�	�!��������4��{�@�u��F,��h��W�s����,ǌ����)!9��kb��`{1.��p�� ��dǇ��bS���yQ��c�7�ɃG߿�qW"c�ݐ{P&���AAU�Ԥ�/�$���� �s�T�?�l�_��41g�aY�y�씄��C"�姫|�� x Uޫ�V��;nh;ifJ���‏^�������u2��*��W��7�f���+�Ze�*�s���@�R
>m$�s�h"�*�1�V�{��V	u4,���v �t�*d�H���hV�=�$�]A4��j����7!u���&��V���=��ج���x���ɚ��xu#}س����F��R�lN4t(� ��ꅨ��H��D��A9�-����X?��W���=C��(�pW��3\�f	b��&�L�ӂ>1�u���t��f���6�P���Zm��ApI2�n�:_�;S�F$A���wZ��y�"���8���c`��0�\�m*/鞜��L��f�� w,K��uܹ�A<@N-�%6���ck��wc)������.p��ѿ0S��Ꮲnn��1�
���g���qi`�ǹ����>�4��ܸ�M'R`ۙ\��l�EH��|]J�e�b�2�~�6��:���Jw�goeܵ�������i�f��-5D9�f���������,K��?5���b�?A*�5"jH�sg��F��j�l������	�.7/&l�����|aU�����4g2�?�T�q~W��Y׿�1X�;����������$�;h�x<R^uY��0PaFrp��4D.��z�IZXЌ��!UQ����Jy�Z��-��$�ߘ��#��	���]+�_v���y{�D29K7س{��vo�d��C��(9�D�!Q�ϟB�RU���,	��)3iZ�ђu���#
��_�w�dؽ��S�0"�M�F�����M��5K*}:)_�vE�e��o���8j���H�04�B憎u���*R��x��͎��"���=ok��%`�����wi �d�Ew	��Q uR4N�����
�����̹�und�']Qʓ �����j��T�r�����^�,a�x�k��LK�!�
m��X#k\�av��#1����DM����������Θ�;(�wx�;���L@[`�)��)w��p�?����ϸ��";���'���f.�^���u�[�t�G��n<�OV���/�������.��Ħ�nܤ������$��K̙O�Dɏ�W�<��#��h�������c�e�� (;��O�P.Zݓ⪟���{!�y�'4,"��U�?�/�!�F8��H.�$Զ���gŌ@/��)��K�K��E�7���u#�B8'�(U�i��pa�a3�&�wJ6bi�
���g>��s3eizH!�N{GRRM�|���M�NW��"B�bΤ��о&�����gU��`��v�ab��5"V<����sN���p�B�T	҆�_���}��C�*ݟ�~R�{(e�<��}<�o����� j����?�X
���0'�����[.
�QV ��1A��x�vH�|L5��_���2������χ�Ѐ2�p��|ClΝ����c�?[E,b#�(�d.+u�L�J�5�7�.��y� ��������p7!�Od�PW��i���\������,�L�!LH���ɤ�1�'��R�����#:2�і���|M��hu�5��}�bG[���m�A��<=+�m�\N!�l}�s<F~!u�Ts.ZԱ��p)崈v?e�_����W7ݙ��F<ƻ�h�ذxGǭHː�A}f{��e��ǹc{��g�j�?xĒ��m�Nk��[��2�C<��9���|6���zYVmuj��C� &?��y|7fc^`v�s��ێ~F�sH$�]G��9�1�YGG*�M=x�1A$\�s'}OT�����H]a��-�s�/�-�mU��*��^����_�����"����4F=���}B-{�\�RL�C�'&(]�Ӗ����<o�.J�9�{b�[�}�E;��TX~|B૯p���L���0Ea��A��n81- 1�*-�Cn���.d5� J,Ww�R��1�X$��]��F|	B�;���Pp�X�m�{Ua.{� ��3��J��Zʥ4$!�ѿ����rg��%i �WS;��[_FAH��̠��� tO���f��})���W�#���x_QK�`J
�!H$��mܦ��>��cM�5��6���k�`ѧu�X��a���Q�����.R,�r�֤^m���]���^g)򋁡]�x���y"��cº��=>��p����r	���><��7�r�á��q�M	7�Q%;֚|w`�+(�V�����3�0���""U���I�Oή�3��s��N������==�xy����̨�۵>=��R�l���o@�;�M�L�#�JyMԽxn�Ab�SC)���ǔm�F�����6����x���1�pg�h�ݨ�.��K}��oָ!�ȓ}���[�b�	�P��Ν	�V�6R�Z?�%�kK��+���$���#y71�rGc�^��D�d�:���sl�x��Qr�͸����אF>���]����u��{[��3�Թ֔��A"6@#|���1E���W+�G�,_ؒ����g�2�1�xC���~��=wT/�����ϫcC��$R͹实�^�p�]laD��~9��m05��� ����/�Я=���F�p��<��xj}q�˵�����(��>jJt87�(�La���%_E?�-NW2,���s�W͛��iQr�4�ȍ�rY��'+�U�v��� ũ���6����������Tz�eW� }zf(��EC���tۡ���"���cL�=�pc5Dh��Q n;�aX���⛾g;Ύ(#�Mh\��t�@ʦ��8�Sj�\�.X4g��Ĉ~�f� �#Vw�rԣ|X�����i��+R��d�T���!v���r|�&R~T"�
F٤���`i|���o�Q�%�ʁa����<���d�S����-���h�����s��}�f��������.���4^@�c���6�o�)P����ٗ�%�S�lQBm�A��*<�e{�-�>�?��r��))X���"�K��-����%Q��2��v;~��r&t_Of&J.��&��f3��n���}ȷ�`=J����E� �#��
HXX��D��;�dT��գP&+M�~�VBq��D0����(�$��
V#d�ZF
֛�l���gꆊa]N��Ap��;9�9�½aK2�.V_�8��������>=/er����K�e#�p�ke|��m�f	_��[H���U�,��4B�����9,�Khuo�ܽl{:66���Tx�CY�	�UJ�f�f2���X'2p�Y1TU��~��eG3G�Wd3$�GHIZ�Oq���`����B���4o0LK�(Fr'Y�t�ܸS1��b��c��?��[A!����l���0l�Χ�}2�C�5�������s<�ZVmVw�`�КcjQ�0C��11�nڅ�y4\ rdzP�%����Y8��}I$	�����D�$:��Λ�rc�H/8�]��e,|��#��]Ѓ.��>��i۷S��/��!R/�o�b6ֺd
A?p^�$�9_UkO8�R����ˤ��]T��Ɖ�7�ҥ.�%�oZ��=�~��-k�{z���LA��h_r��Ay<O�)��|�z�JJa�5�<6x�c�G;N;�d�}�gkfbɉ6�ߩFYQ���s�Nb(b囹��F�p�<(U8Q�i��>��N�'�����G,�"��͌~
W�ף���mD���S5��!���IE�zò$D�	u�i=G^$�fY�.�$,��(��9�D��J_�wR��g�m�)S4x'~����9�b�1�i���G��Ks�P�4�+�@�c�]X�tŌ��Hᨓ`OZ��""����%V�mH%cL�� қ>LU��ih�.�Nr�Y�|�	����<���F�gT�K%^X�'�gWH!�ڬS�&Rnփ�̂ԔZ���#��aQV3gA���9$���~���Л�.�,z�%�*Q�zS����/`@2�*�}/��̺~��g�׀�*N�u��{�Op�B+G��{��>\ҿ��ס��)��4,ǭ8�=�JoS�o-?�̘�z�W�oj����ͥB����{�ᛶ
0�Wk(~n�k�u�Y-�����%1Q|0>4� ���e����F�^(v�mn�V�����dŦ������r=Z��']ܣ�Ú�#�!�\4TЎ�vN~\�C�,]���W���]���ԭ
�h��[|�\�N�غ|����0� �&�e�ŴKT�=7�J�=Z-��J���WU�ڀ!Y:�fV�\��\�+5*��zp�r7�M��T=�P�-,]�(k?g��ם�ŕ3PFס1ڐ�-�SA�q=�u%H�6v�}�9�9�m_�%{�M�_H��&пBĶ��§�r�]M�A�(u����H��o����eϪ�X�!b�N��&����^Nᷞ��U�yj���R%�>\�������]kb���=J��`t�@�>7yʆ=+'�[����A����j�_P����$]R�*|NN��N+�|fi�ÈC��:΅��
s��"��a�-�-�^��G/$��-r(a**�jT�l��KP�V����T�*)�4#':#i���jp<�ۂq�of�e���f��膺p��a�ƞ�Հ%�R�58�p���[��R�<f%5�E�[�EPT��]�ܣ{�	m|�5�FLS:����X���Y��%���G%T�ؿ8��jz�dVwp�r? ��z_�IZ,jʞD�gfu�_�Ο��r�$��×{������ϩW37�%hj�A���n�?�r�F�*2%�«ߘoJ�^,r~_�y������d��d��j�m0�Oz-;�LK�s��������)��y6�oڋ���H�,�Y��/����c�;���V#��m�.w�q>�y��";<��y�pʜa.��� ��.��[�k�=�}��=$4 '��/�P��Uܣ������J�*v��]��2v�"���b]7�#a4��a
��H����ҍ���m��C�R0l7G n�-�&��M~ ���\�¬R���Ou�dTBoN���S�#~�
x��j�h�,|Pŉf	?�	J#l^�0xk�D!Wy��>�[s��$�r�M�·�@�.;!�&�Q�=�]�-��jY1i��v�a�)���?����Y p)�e���WI��=��[2U|6eP�4��ʈ��dc �*����-�T>|�Q��!��l���B`�f��A��>��/�}��c����]���``i`�D��1��@����@(�G0*J�!ʚhu7��c����}�\���Z'�z�]�⽚V���?i����/�oe���0��g�����4�`@i�ѵj�bP:%(T������L1�4S@���\��?o�&O-��Bo*X�"!Ul����&��u�M��(L��~UFXܯ5T+�.���=�#�� ��u ޞ)�(Ty�ْ�g��G�����c|(nan'!�� I59�Өr����^Yf��`�K���u�n�u;�R�$��YR<�؀Jz�+g6=]�K��P�b}96��[�
��i��UE�B��Q.�a��6�a����>�,��I�4�Bm�E�"�6�9�Ό����t�ex�z�����v�c�⿯/� ��]T��Zu��Qcp3�[�(�o�L0=T������#"�`�%��	� 1�U2��r�+��L�h5$�� i��Rn �m��|V\f�|a�j��"d����v!tX�V�l��K�=�n�C ?ȵK�'T���z7�?#��P�h"�m��`:�/0]~�m�D������&��z�N���<���G�-D�2�l^�|^@�|��f/�F�C�Ǟ�C�_�-U��s�ԙ��͈]Zx�;h^����c��#�$�7��쿔W�ǭy
����@�̧K���%�{)���xL�-��{hp���wYڠ5Qא��=�n�o%0!$_`�]61	@8�=���3�m����g�Bw�v�>c�|��U�N�
����/ L�6��>�Æ�-�G���}�c����)���Q�S[ˢp���5|��n��/Y�'V&y\�\��QCAm*dU�!�R���)��o���/�5�Zzbж%x��b�� ��F�8����[��qv�	�8Mr s�-䏙T����	��5�_!��33�pT/;�Y�T�5����(��=�wȳ�H��t�\6�f>�燚�Gw@�o�zDZ`.�y�U33:��?�L ����,��P7�B�O��z���V�l�6��	�'��^w�R����*�c�ɓ !@��q�����|�P���5�D\`���P ��������N�}s��9�#F��sh�5mK������B��\,��9�-Z�{*��D�E�t�%�x�5���MƵ4E�X� �Ԛ��*�3u��z̯5�#�N�j�&f����S͌�NR&��60��X�^/�#�$z9�b_[�\"T#N�_�%5 ��c������LT+�3�p2��ؼ>{]�/��k�e�D;@�V�ZM/�"��~�����tWd%s�R�yu-��du�`W�寠%O���͚���%�-��j&DX��f0쀹�؈��I� }]�v�)I��	�G��}����]b�J������G�0Y����E��ŹU�0���L��뽯I鱒�t$�6zk1�o�_$l�޿�O�\��*�.��|	��:[%�BOz|n�ɻ����d�="���Xo��y�}�m��g�P�-Wo>��Yj���'BZ��M5���PS�sO��Z%�Ã~.��X~�s@D:��y���Sz~�ȞS�Y�3�MFe���d��`��,]lƍTH��IwKx}�G������"�:���Wo�Cr��m�] ���+�K%L�p�w���+����
�z�u[��F�i�亢��\R�a{l8���ᦦ�xQ����E��\tF�GhN��?����p�C7�Br�`��,���^Q����k.�g�Û7�2�؝|�گ�߷�͗���#W!�aK�鹸����޷1�N���G_��q��`5#"�3��lל��}����_@g��9�+zs��ۂQ]��M��a�߶~�^�z��l�UR����7�^�ޠ�ߗ�I0vZ����S�Il�N��Ja��R2<@<o�{�s�feH�(��U� k�]x�rs��,z�[ ��Fֺ���)��̰��ozrC�{Dن]�p�N�0��U��|qX��gMu�9��RN@X�B9���	>�&6C��Ģ9Ǎ���^i��Rcm \���]X8�[�..�m���\�R'�%,⤗���C �i�ɑ�7��=�T^�q�_8� K�� �F�>�um*ě��dYG���Y�&~|==�x�ܐ��Y���4�ٝD=e���֧G�?���V��X�b�S���K��������y�i�1���7���x�(�N?GnW`eKn��!�mpJ���|�@�ȍ2�'�,u���&�l�|8�[V#��ctW�:�Ud�.fZ� ��K�� 2�1�����ei�L.�W�p`:H��tW�K~�}|:����T$�Q�JB̸]�t�9_Αd��^�T,�r���"�XS��dn wm7`���(�W���g�C�i�-F;�C:���D{m��C��7|f���^	�L�L�D1.]3X_���Y�ό.uY���(,'���W�;�� �wLG30�Z`���鿲"��!��e���T&�E���R��;�a],�O�t��BA��>�Y��]Z-�J,��J"�����Z?v`$����iX���3�h�e��y^�4i+��Y1�  ����K�oA��	��<��_����ſf3�Bq����i���z���o��j�j�x"��u"dJޗ�aV�8aJ���Į��![(�B�r���4�o��Nq���1)(��X��'W�����X+˾m����DD�)�!�,�,��}2�=��zؾc1�Z$���#�q�V0~I���3�_�eW��HRQ�>��O�\�W�6!?[l
=���?�-�(�s�~*��%/��}I#ug<XDx�z�#Z7g����)�sid�9��lL��0?�/g~�j}v>~޷�k��U��2�!�a�I���xRiH��0x���N"��9�?�#�}'�K���:m�`,�z1Yh��H^̧�$n�t�m�����5?�-���l��̻ZuDF���zr^�Wܙ{�1������b�pRMNJ1�B(]l�I�H����"+l�4�e�!FsWq}'��F�uWn]&�d����Y<�,�����p0#,W�M5�WkkQmw��סA��/�h�B�*[�jὰ�˃b ����+~~�-b��[=��ur4wm������b�'�2��!��e�����W&s�B�3q���E��q=�@,���!@�>".���a���!���Ι|l\s�ƭ�M1i7�A�#����
+�f��5����Zv&",����?R[�<F����,��;�7�7���#��5�S�W�3O��4�W�����Ƭf�j���9Q�w@�+�Y2]���;v�V�|�Z�����c/\a����9���_]��flyj�D�}&���'`A��W�j�ïE���ü�F�a?�y(<�ƜX+�z]��^��5�0�����g���L%G��)��v�UV�$,�]��%n�X�����W�!=��$����.ƕ�Id�f���4(RWI�dXȬ���׸a�eP�QQ3�\=IȬ.0�g���-ߤ,��9��\��5��҅r"4��`�lPy�_�P���͍�b�|@�jJ[�C��d�L���?������	����b���m�z} 6�r��Du_E\��2��q���������?��f?�A����A���0�pJ��O��KEdz�x�y��������3'���b���ï�)���i�국���D�>�T�e�Q�&կi !�����M{ �4�D�b�jِM�^�-��haR�!��ۅ'�1�
�Ԑ��4�;0�&Mq-���E�ku�!B5a(�7|ͮ~ -PAwq��	=a]�VЦ��I_�rE��hb���	�Ҳl�E*m�B��92�x-��J�L���4.����9�	�(����,$�ko�u�d� ��1؅Ƿ���'ٮ��=)��↽B��%!"�;V�;�Q���?."���+:최��R@ �G=�
'�hq�S��@W?v�1�D���S6{�K2mb��83�Ǵ��Y�qÎ��CB���� Q�;�#Ӣ5�k�i����S�s��~q{�`�����<�� 0�/�e��ʾ}��!��������k���W@��Ik��>�BC!sz��i�Sʖ�	g>�_To*��s��5�Ō0eN�C`P�����s�4��� I��OB�p�2vV��i��R�,�#����F￟��`,L��w6~�d�+�觺@J�|��i�=��[(�	Q�F43�'�?0迈�<m|$�N�t�z��TR�n�� �z��ƐTu,��忒�vz�bk%}��B�0r�9�d��}$6��j@����]ۗw&~��o��Š�"�}a���!��$���RK���PCk��E2א�Ln�p.q	�,��#��򖞏~ k����5�J"	�~�`5h�K'	&P��.K2�( <q�o�2���3��!�T����y{O X�'����|YV�R4B�✆�]�F���_�LcSջ��AB
�BqA=�?,/-���Iah$�n)���9�x����3�'4�c��cZ��a��H��|�8��f�i	�һ�2���w_�
�e�����u�%��9ak�� >�u}���F�>�C{cc靍nsi^6�I�$ϕ?Lf���7�$�iCϻ��L�j��tm�Q��V:�<<E��8eo���#�=&H�4��/F-�Q�y��Sa'1>��+��ꯠ��KK��F�V)B|���ʧ�a{��m�]�ؓ�ʹ�������������EA3���7�� �TT�̈́q��T��=W�K�D.~5�V�(8���M2�$J���4r�c^�Sє��u0��^5W3��L��bw�a�.ԅ=Fڲ�I��8���S��*wW%�n�BO*=��}GIA#P��m��+]��ݑ6��r�sC/����u}��.q���zW��9�.��:�Y��T���x9C*�:�<�IH�Z��2ME��cvE�Rm|r�U�l8��m8���ҩǑ,�I�Rάi��OWmA��'�+���0���=kc���qK'/�1�U
$w;S�e�� Y�B���v3n0C5cɅ����O9��@�1���|T�۳���4xA�A�+��Ǧ�ޗ�<��~���m�Ԏ�!H��K����:0#��;�J���Z�N�g���� g�s����߂�7c'�2�r������Ur��ʳ�]�R�����$��kz�vM���N� ��yK8�8E[􃣷���7k�����p��Z�T[4�	�y��DP� u��	Y;�J%sm��`��n�0�l�m%��$�/&�P����E+��~d�I�Ӕ�4� �\�:u,&?)v,���W{g̞�A9�X�p�A����5�r�8���55�_�._:@�BYShSo��xl�%��6ɨb�������yaW�뫶��ҿ���Yno٩/�w`L�=o����׫��5�ʇf��G��j�hW���=7�u|K��<�;]��T��P&F��B��q���Ӫ�E�u�.�����=�����}4�-��Z�B�:���ȹ���:� �4�gEb��'ȏt=ۼD��y��i~���U����`�
����y���>i�iG<m��LGICY��o]���_#'쁐]A�6�������H� ���%��/o�����k-�T�𥟱w���[mT|r�����{��~�A�8���.��[x�
����Z�&�I	�n>{��љ�z˪k�i'� ��7|��?kߣq����UR��ș���� ��E
!�"C�h�U�o�ħ3 /�L����s�m�Ȑ@��2d���ӎ��<F�巽�}�����u@�����a(6�q�g���o/
](�4�72��K0�+Y����jK1m��ږ��&ͺ$���^�����in��b�Yr
�ＪN^���:@ukM�BKa�q���ǜ�{�γt��JoѦ�|�s���������*;�<"�X�}E����tWf�j�cqݯ�S�p`j��],�6��-�ڊ�!E�"f�`cT�x40�7��������_f#��R�;�f����\�C�����cƿs�\�(�Q mԽgc�ْ�mL%����s8Em��I.���^p�)M�<�0U!04qߣh �哄&ޢa�kM��#���0�y�[ૼ>c�+��~�G]ӵ�5_"D-�=�>��8�֠��
�u��S���%�ҭi or�2L|��H��Y��H���6onU"s�f����h��b��&�0?R��K���<���,������}�>�;|]`����N��*�s�Y|�k�=bn"��e������kKX�C�0��3��ԱC6�w�DȤz<sw�w��^����s;\~�3t|��h��D���r��8����H>y������d6?��@�h���k(����?s��q������1��z��z���%�|]=�!kR�nPuE���'��[�z����Ǌ�n���&	��D>���22A��y�W�ACXiO,R�s���g��'�dŰ:��6K��d���p#{�7��#[�D2+���!=����"dU�WL���|���h��^<K����XN�3'l���i�i� ����S4z�<p0:&�]��I �����K	�BS�q亖M���Uk��`8X��0�"p�8�-
fS��@w#��`���`U�$����`�f�p���<�zpE0�d7�Fr�r:J^���m��[�n�)>��b������ h-~h��=S�����aVm�?���s.��Vz�朅Bf�R�+��aK�R~ex�<b�3b����a�2�r��q�h�3��8_�����k:�������%�t �#)i�Pᄬ�F�W�nt�׷���>����p�5իK�.�6"��:�E������"Z~�Av� uϏg1ݎ��	3�n���o�`��G�00�m��ї���k����� "e����'i��8�wj;��ک���6[�K����x���#�H��*���kJ�4E���&���)]t:f%�|�Oj�t |�>) 2�GA6����|��)>�{��.I�8,��v��[�v"���/f�d	sUk���4V%�t����J�Ub�c���k�@U�Y$)��r���ҁh��:�Z����꟤�*`�rh4�.N�~h�I��C	&��0���(��}��Za�t(]^���ӻ�h���tQ���u=Gwƙ+u&m.���ΐq�H�-K�{�~k�����8�R�7��4��?ag�B��:���`�����3�Bb���u	���M�w��I�6e9�?��.%�J�����=��sg�o{�^63����4ϟ��ԯm.���u|D�
0�tM|��u�YyY�q�v!��B��	�G���7R����u�"J�Qj��g&�./6s?��^��%4��V/;��*6�O����%C0/��-�ޔ@�&��%Y���袹�����
���:��{9>k-w�}����U�Ŏ~�30��K�Y3����6WB"On��<��T�У'-Qt� �A�W�s1�%&�q�Iے(5&��{#{▆ej��Y����a�CY�K?��f��yL������p�zʛq鎝(� [O��^c�AD�,Ŋ�h�Pq�I��sBf��o0�C)�*8'(�K�o� �i�F���
*g!<n8�	7�D���s  ��6؜�ٶu�E�6)��7���L�~I��!#e�&2���ܺg��$egL�Y�4aH��=��3`��v	�>��CU���ce!$���ԙ����0kϨ���4p��+s����}y�6^�/C��E��(�X,6�,��,���$� ��Y1+���?��Y�&x1R*�~,�a��a)�/�:��/��,��Dr,�p�'��qO�K�p,?�����iSd��'�S�Jͩ��k�#���_��{�l��d|P��c��Y\χ�|7�)^@���D����"��X���;��$��A�\L��'	�Jˮ2A�:�m�7>�:+�V�4���ǥ�˶%)]	_3���
��IxY�R�*}r����#�;Cק�B������j�)M�L�Gʿ�R7�0�휙:�ܕù\%�M�p(���Մ` �;`��?&o�Y�p�gD�쉥�Egp
��+e]�$��n��"T��� �	��d�A�s���Q��!(�_@g�ߴ��+�^�:�~�`|��?[b�!���>����3��"S](��.��hSV�3�Ɏl�u�
��`obt�a�D���M�ii��Q��b���Pfq���Log6�g%��)�i�"�>�H	-�޻��o�$=��AkÉ@��d���F14,��s��D���~r����!���1*��LF��,H�9��3�w���rb;/fk�f{_a��SU.�p/G12ݱ
�EhV���U�-IT�W�{�ÞD
���A��3/�D�҄q(B'��ڐ���R_� O���U��w(�rx���|���S����N��/�eF7�T i��=М�{�JǛ�D��.�� ���`�A�q��Fm�n���}�)�G�ҕ��,��r�)��$!�l˱O����2Ag�F��:�+�_�=OE���P�Stg��O��f�2���T"(zC
E�0퍐���Ƨ�Bj-�n��?G]9Yuԕ��/`�����	�:Z�5����Y;�S��z1��'�Ŕ�!87�*V��0u��"la�����M3(����x��M\���ҧe?�暦$Rb�v+Ӊp�:�)��<�*�g�=����
�8�e� T�iq�?x	{?�;9�E��t���}7�"ՠ3Ka��P��0��sǶ�:%�"�B�	C�W�2��T�Ѣ�F��ʲ�Q��� 	>�}h�ʳ2�Eezt�b��j��ו�W��mB֜��-m�<X����c2t5@
��&j��fY�Ўq��2�bN�5�u���Ĩn=|����V+�P/���Ľ�r�d%ikED�U�F��k_�:@!�A�S��1�&�)t�5�8.�F�|����u�k�p 0 ��v�!���{�"�s��@vx,x�]	C|9��G�Ǥ��.�'R͔�8Ifh�)�?2!��13wJ#�=�qQ�@�k
��f]e�p���Y,̵T�W5Q��跘"�8���K��3�u����.l���.�W�<�D�^��=�"�xz2ަ�L��#ob�m?Bs}mFf�ZG��h�F�����c��ik�0@�~K��:��f����;7�t=D�b��K�w\���Ѓ�_EuɆc��>���47H�в��e�F�*V�ܷ�=g��9�h�ҽR�Hko(5t������������tk_ɽ�&j{��ר @�G"��$�m;��15 �a���ޤ�0�B�繳8E]��̣�3�"ﺛ��zt1/�����4['@���d�/|�`am�#[s ��d����9@���ں:0�h�j�4?j���F�8';0�|����F�D���`�����'d{6$*1�^��X��9�"H�+C�ڶX+d@������� �L%����"j�
���� s里 �vk>�،�k&Mro�)��z�ԛ�|��oB����G9pbgo"�1)kŉ�J�b&��Y�d�ڜ��N���R@3��ܴ]p�*Қ-��ӄ�w�^q^ل�Ea�P��V)��mM���!gb�,I�r� P�<+!���ވQ�Җ_A���F�tBa�D������O��vV�������%�m�I� �р��
0�N[N���H��Ep9�Z2��1�ｴ�Ot�j4I����0�,��JЈ�g�l�66Y$�~�����Ɣ	���ە��g��w�\�����e�Z3�2��t������*�8���*W���M�����VU��r��a gQ��e�e,ͯYumڭh�Ӷ��ԫ.�&z�n�-�Kҳ�_��`�bL r����nX.�� nm�B^,�y����1qn��G�Ļ�+-�뷦� o�A3�O�hj�� n�y[��T��{E��@����@EH8����M����I�ڜC�i/��U��y_鼘���2��n��{H6���Ѡ�:�
��9�KH7m�/-�T?�h�+�=RU��E���偱�	��uD�J>~�l�獙�H��\)���1D���Yw1�R�bjw2Fq,ɨ�ޥy�p��M&׀�B+��)�K;�`��3�WI(t'����A�B�1.�<_G$i���4����.�*�h>�J�vN�uݽ:+��#�F2���uE���V�b�\r�ƽ����7,[�_�ї�I����P�ۤ�>�`��ڴٿ؍h/CF�"u3&#U������r�
4�?��n�^{o
��7y��a1��Z�J6=�?̄xx�DE��78��V�7t�^���^k��î����� ����yėp���5%zG�N�w��'�~ŕ�s\D:m@8��-_l��D�S�lp*F�l{��4��vk0����-}�oҦ;<´�eߥy�����
c�Dzo��l��ڋ¼U�2�����rpE��F����b%_`o��`+B���q���F�^���	韻L2Y�41�*����8�P<hL�z��oCX�:�!%��T7�+��D֐��^�n�*���xIM�HG�5 äC��V��x7&�BHu���D1�S]<�s���Ō��V�*�d�
���N��2�v��,��>�N�eK_��Ms�Y�_3|��� x�o��J��%���U)V����@�z��{Z9�RD�z}ðOUW����d�cb�=7��e�\'�ےR��0i�\.�\�з0MU]��)D���a��4<�+�GM�Fa�L���֮yK�����7��[���f>�v�Z���B/;��ݣź����@Q�p?�]�y�����>�/*~��z�ͬ$�|N�N���#7Ҟlq�j0�m�٥$>Y��!�zb�+c��T���8a�C?�;����NՓ'B��B�7�����,�l����`v����h�Z}���\�����[��������O(wwB8� �e��6xۗ�����
ި�p΃q1jA����QX����z��I/�#o�����uY����C���+��K����YIX�RZ���CA��n�V�	��2���69�˄b�x_�@�Љ�_��K%�>(�(Ϸ�Q��m`��ĎZ�_�q\�;�hp#!�>���ns��񤲹E���o��Q`��q}����Բ�4��7�h�x
cf`�������7��r��L-C�҉X��ͦ8�1(�ĀHr��)���&������;�.����"&�̼/4�*��3�������J�sB�$����s =�+��	nA�F"Vb�2������I���z��N_&V�����������؂�@)�θL�(�������損�%��hua��k}!��&��~zie,�'�+.�v����れz�P=I�����4�%@G NqR>��~���y�oq�����&�=!v=���"n�>{ 8�{�eJҨ� ��͇�c�U�/�f�e�G��8�V�Z��a(���'m!�^��{˕Z"Q�-��hAX� CJ^j�9��3 ��J�B�A�t���2�v�!�9%^�¹M��S���P'P9����?��f2����!�����	Y���xV󧾣Cʈ�ށ'��򤈳��O��`q�.yJ��i>�Ԇ}R(ɦ�I��h�D���b��s	A>8��]�M��Y	O����HF(��M)	ա�%�%�-i��!��j�W͹���,�� ���b`B��V�֏ɱݡ?�N'�+�-�0��m�,��K{f��YT��dN�/���%�,xX�O�i��@�sA:HV��qG,$�j��!��	BQ�!�W���㠫e�m�I+|Y�6�����!h�B��`cD�Q@j/=�n����my},����_�n�ٕ+?d8�O����mec|x��nш_Ւ���ӹ��B]9�8���o/��\o�O;$z�*E����*���up�aB/�؛�K�:vB�h��\=���^Y���1���4����*f�E[�8(�T%�%��M��w�H���Z������7 � �EM��#R7N/╮(S{��D�Z	��࿌{��W!��c���G�B�FUcy$ې十BT�Sx���|cY�c��;K�I��_�ց*9����e��xy@K��=���ez`�Q稈+p�vcɴՔ�S��R�|E�Ɉ��!	��Csf.Oj�HuY!�p��7vM	 =�_/����bt��ufX��̲����$��v���^��ݑN��3S�����^��w����v[�b╕�ƞ[V�HsǛ�p�F���ikQ�� �e	T�
��\����#� A�r����@�8��}T·e���rJVN�0��O����A�5Ue�'B���A���c�2������r�lYs����ʈ�D��{�����b'e1�Ch���6��C��0�Gɞ:%�7��Խ�T^��Yꤕ��2�$�L:;N����r���d�P���3 �z9B�(K'G�1���L��k/�m��w�¯+�)�G�ő��ݓI��u�až��ګ$��n�/-�^�C��}��`BxH?��b���h����@�j��;���>hc�1��ާ0��+
�{����B�f��.Щf��}��Y� �F@!uSK9tR?w�_�}�<g�Y��:�z�j[^ݯ�$N�K8�B�$4e��7Q�1\�K��_�*�T9�'�{LSc?_c�S-��b�H������P䇬���@���P`u3�EVT�Tb,k�_ݥe��p��t=���W�$�j�+g�;�@�9�2	z@{��p-�bbM�Qj��0�g��a[`�F���/��$۪�6x��M�ח�aD�b�i㊋��^Q������P1E�U�Oi��vB^7���X�TB1�r�t3�&��S�Y�s���d���o�z�9a)^��]8�e'���@gi�\�����/��h�.��e�y�n"��71Ԉ�I���z=�@`
�P�T���i�N��%%*�m!�h��d�-��
��fO`�:F� ��Tetq�ߨ��dH��Cբ�����%Z����i>Z���_JQ��x	E[ �z�L��e\��+�/���E�3R^�$#pE�������*�3��k�9��-����Aբ�E,��o��cy��eW8|�]��R���;��t0�~N�첂�;J��b�rV�X"�q�����H�Ȇ�:�L� �E[$�MOuz��d�����zV��x�k"��r�n[p@*y�6��XkG߄��!���a�e}p���X�ڬ��:���j j� ���B�ֶ�A����kC�']N�y��o*�����0�ܻ"x}TL�O_$ Z�X��պP�&���>���c��HSH�|0���W�q����rTj8I�����'���F;ni!�I{|�`ַv�휧KN7��Y&�';JsV��'�?rF�_HW�&z�M�v��ס���d��Q<�%J�%ޣ-�n4v�m�[Ϗ�"�mʹ��F�Wj?>b��|]�mm��[��x��@�U5H�YXP��6�Ķu��|��I�%�R��?�9��uK�k���)�Na�!� k@���"�)�����&�g�Dk�H�/��L�+W,qL=��#'�7ʑ'�C��h}��7;c�N�DF}U�v�B��WA�]�/�x���fe����2��r?�j���sT~	g�M������2�:��V�q.Iө��4��sf͕8�nEV폫�6���o^M]&�D~wj� ��$�BZ�p�X��`-N3W�ф��Z%���S�6�(������4�[���)���1Jc�j�,S�MEJ�����g�� ��mI��ɣq-#V0��;J�yO>P�� ��6����F�B.�W~�� �ٹ��.	��$[�H�&�g�dtkv�)�%�$ט�W�~V(��2ף��;�Oe� Z~Sݸ@���&��R"��Gџ�3�idG7Ar]a��;�LNuƾ6h5�i��Ty�O�n�������6�է��]/�V���<݄v7�|�0�g1 w�b�z��E[&Py=XgV���Q  ��<�u�-u->�V�%�:�Za�-���a����N�Èi���gb �y�@�↱;�P�t����s
�o��L�a�`o�t� ;D�c��o��zM_s���LSh�Pu�,W��1QJ?M������F��3z&&�6��P��������g���	�+�]+u�CT�Ζ�G��f���utR�X�7�tS�	�T�SwW����s4��Y�+� Og.n'��+��C�^5�0�� ��I��^uP�W��p�1X�'i���Y~��f����\�Q���vj��^���M�8s�*�U�w�*��0��K~��L> ű�i��)&�A�����WaE���s�9�h�J���0�{�����ՔЙU[r\g`�/��3�'DV���q=4ſ�A{����cϤ/:���V��:�bѷ �����-*ٿ��/]�w�d�4b�fH�cXWj��+�v��ǳ~~Y�>�� �$g����bǕd���n��zo-u��\���Ǝ�<#����o��s)E�W�T�7"	��s��%ȧV�v0�g��`����h�/h{#�H����i+�l��?��$D��Uo�� i������s$~��ip��fG�k��5H����ť9]�wW���/�[�f}�+�k�$�*�e�0����A�KP�C�g�O�o�$@`��2I>n*0p�)`�����u,N�(�$�3��ե̜�ͪV%���M��R_�򃼁��('u�Zm�/�苐禮�1�(�����ȉ#��w���Y	���Gy�W�3
��{"�BWiR�?)#�
���R�"�4e���
ʆ�!�?�o�޽[���]]��/�*$N�u�2�>�E	�麺rh1xǚ��I+��^ $_�L(Z�ʹܝ��v*���$�	^m?�\�8�~C\��F�tؔ��+[1|�r�O�Tg�]ƞ�!w�&פ��Kwn����J�zҴ)Z�	��1�9��W�m��Wru����1q�4�Z��B��I�{�tuT&0j=���B|�d��'!��*;1͗+1m��sq�[�k^:�ly�v4�A���v�f4%��A��S5�]�'��=�E� �S��4	�]�X���3�j�f���p0����_� �L�w,���d�m��J��E��_�k|X�"X�Z��=�]��檻�K �4�#�6{ D!�E���[�ϸ+0�HJ1��/˾�x3��)�fFiT���8� �]�Rئ �H�s�x�dTŃŀ�v>42����v��c� ,�:�Ser�5�`O�i��&:H$h|�>%s����%j�ٵ�~8H�RC�2�2�k/�q���xt0���aUݱ%)���,:4�fǇ����.�	k4���z �tW��sO�Og�m˱yOP�rTı؎�����t^�An�Dy�߭��8l7��H�;����.6p���4�2�'A��㌲zX��ڧQ��T�|�������C���w����Q��rb[�D�s�?�\?� CG�	akI�cnv4��B�}.��@% <�8C8?.;c�qޢK,�@�?w�C���lDu��|mgW��� w�U=��\�%6�^��0�.�lv�Έ/�fY��)W�*౮��
�ϗp��7���ƈ�;���;���K��Y��us� g��!q��\���v@�� �#̩�l�q�6�(�N|���H��[��-{���N�
����r�:uS�q��q!���|��6���ƺB�~mS�����z]d�c`R:^Nr�-�7X�ʔg����ա�7 ����f���Ϳ���y�oOW��kL��C�D��K!x}Ȝ�E��PlH{��=��av'�X�4�J粏v7�r�	�)4x�������Y1n�*tZ���l�?����f5ǆP3Q��4��|j=Aatyf�{@�Z*���_��Wh�zp���F�a��3k�Bu�7im����0z�򪆞l�?�����6]1���E��dH���H~������_���t\f�����*�r5 �غ��l�c~?r�`��cY�ݷb���%읃�D1be�\n&�&<��=x�r^�2m}{�������3�=CH+�G�\��rP�Q��+j,țW4,�ۑ����:��bGQ�	{��n���;L���A����"�k�Ð.]�\E>A�g�q��6,�X�^2:H��	����3n
/�R�@f�9-���,f��"�߸4� �A/��268��1�$�mn�j?)��hS[m .�e}�K����A%?�����2=�V���*�-w0	�7�ۼlsȃމE#�x3R��v��w	p��4�����!g�U�'t؎�N-�GɎ�B������kE�LD�6������1藣W�7�0���Y��y��g7�z3�QK�8e��#�3�i��>��?��A��oD�{��/g鑕2�r
��ģD �LМ��|Ӄ���]���]�)E�$ ��Cun$�g�3�}0�>g�Ԯ���+�]'��i���?�����k6qM���3��uz+����y�29��t�*B.��^ꝏ�Î"�P6�����WT��5������;|�G kM�\�� A����T�=�T��⪴�*N_i�lԄP޴���͇�b�*gn���7U���Я̈ �臩,���bR��uIm/ ZK����MvV���A�4 s6����*4�)M��T���1/,���i�6u�`��_����~�/ʅ�n���19i���Y:��Sq1/ZSKtI���c�pРIDTY",\:J ����(����N�i�em�}�տ�8ig����gf�ъ�t4$q5ނxE4�:!�]���e	��z�K5R��ܻ�FTO�
.�"A��];r�m�)�p���"��.��QGoq�Ľ�x�����v���Fy4����ɉ��P��;�k����q_vGw�e�@,�f�4��G|-OR�<��+�k�r�1ʈ<Df�L���CZZ�MLy�0KJ<+~*�ڻד�Y�u�q%G(��wY������ ��L�W����SN�W{�W��胷��J%Z�O�\���'�·t�S�yK�%��5�r��C?��B�%A�p$�"NG�����rWH~�셝��
|f휰� ��J�zݴ�[��&$����j�S���O�Z�'�9�� >8�RB��}��Ц��������O�r�.����|\���
�����JU��$M�L�(�L�3�O	"�y@>#��� ��
��CVI��ɤ��\� �J����Хbl�6A��!B 㪸E5e	����E)���9�s����3zp	3�����5���I_/�}B�wc��//3���3ϸ(ڎ��>�����H �����0���Z����d�;�B?�&���Y�	A����{]������?�#|&N)����ղ���1a\l��=_��QB�1u�'X��2�@�-�(�����2n]o�v[�D����cn�k$�y�}O��\c��,���Z�k<�G���C?�B$�R��sȰ�
S/g���2��-�q�B�Fv`��E^J�5G�B���b3K�N��iu�n�^@| �NDC��Ne�z����O9V��dQZ�5$TVf��¦w���>BeF��E�E\[�%C���6B��妴R����a O@�%�1�9�8~�W�S�O�8�J�jU���K�>��[�v��rӗ�|�XC)ҍRI_�B5b ���J&��~�Y]�N�Yp�q��Ѥ@��d��5Ĝ�;[$n����d*.�W�g�_�':��>H�3d���t�a�*��Lں�h\Vx�d�[gȦWxO�{�����O(�NQw_�C�b`�|F1��>��'��Q4=�x?K�[t� /��;��;9ki�����;'f���x3�ޫ���f<�3|yCJQ0��e�"$�@F����p��)[��F3�C�㠆�?>&,�撅��T�lN�W�����.�cFU����_���dl�7��@���} �;�����G�C�Mp"h�[A{���;0�@7L+&@��q�f�9
P���k��[3��K�Sc�_R��� �$$@��^)�.��*�����;suU��6��T�;e�f�L��px�ZT�3��A�yL�av��^V�?�{�$�|�%�>Bl���fZ4㜳1����L?p����{p-,����������u=����ؓGLM�~��9i�Q,�W�j"��ա��f��8Υ��B��YY�]a �����J^v����L,t�@��Oh���:"+��ui`X���������������>��߈pM��"VL�@S#d߹�~+.��2�>>���.��l�n��jǶ_��6G��S��ELDF1C�Y�v{Ʃ��2������(}3�k�@mOuk`{�W�kBJ	���� j ��X]��c�x�����&J�h�tF�*:�
.T�u~^9���=$wvl��V?��\_�Bi��"@��Zq����`P�H�<6�E;JM@�fS]R.���f��%h�J� n��
��*����{+���.6𛨓~O3S@��O�gn~�G����y�/��f�0���5^Ĺ��ɹ���H�}83����mKHb��'�<�u�F�d�!;}������pﵬ�
?3����u�k�͋R\�@�8�f�!��̞�R�q=�LsR��ٚt�̢�
�����C�Fb$�R6M�������9
�E}n��v�0��~r����:�q��?*�G���u����Sj�P�!��^�^��)4�`�*pf�`ORB�q�����;m�/ ���E:w�l�=뾎6�p����8D��?��Q��?�O�-o/�L/�")��ٔk�AoN�m������f|F���� 6��9�I�7͚* Ɏ\��pǃ��n��X�l ��L��p��>��}�~�y�����A R~$�1*�6|� R����z�����_�����k��W�s�xB�^}I�}�C)p��Y���_*ؤ���W{�6I�Qo����`w:M<�d{
��J��]W؎���@LH�SY��4�-����,͓���SR�M����G������X���j{ eb;��VrE��uζ��to���s�W;n9��L6a����N�qO�T3�&�ca��2vcj�K��ߩ��̼��	���A	�}�6s;	�b��v[�O(ϫ!�7֝�z�xuhoR|p*#��y(bQ$�?���*���Cc��b6B����,8��?ȳc󷕥/�i�E��{�رk=D�h-�}�_��ze�_1�\��&�q�$'� 2AE��8Ú"/4�#��3��g�u�Q�#�S-���g(�V��_~(�i��*��q���F��*ٞ#�Ff���u=̤�m=I�#����盉��/fЧ��Xr,7;Ň!�|�o��5YiR��=\b�<~g#�uӻ�w�⊊Y����z����?��۸QDI��fU���"� j=[4o��Y$��dwSF;�K.��T���Z�\���� àd�4)��:���Kn�u�����b�>�6?�^K�P���n�
!mk��3N|� ��.^����!y���xXX)����3l�l��CT	�9����.M/CA��Z!�Җ��3̥��u�;~��H1�	���,�a�o��+���O�dTX�{MB2B6��af�<V��t���,�����N����������UD�" ��X��+g�ܯ�
(HmKO޷w�p���3{�e2��2���4m=��Uu�'�Y����&�`���
��F}��c���\C���n��o�#��,��-o����Z��	\Il��`�H�#�4���1t�l��W�S���9��~��5��+H�
�LB�g�){K��P�GLFP���p ��*M��2ҹ����=�u���Bi��$ʄ:�z"c�������m'���]��V�vk��o ��"�h�^��T2���1_ɰЪ�d�����)^�ʼ�Y�-'��]�"uw��I�qP:A-w�l���� R�,j��]��䋊GL�!��ހ�c���g�a�#��;�~4��ؙ:��Φ^F!R�-�ޟ��?$u]�?6%��>�]��� r��~>x��Y�k�6.�����(��-Ҡ_z��k?�ZxR���2՚���AvR� �mQ����m?�7V0��%�gR�ZG����>����IjQ��T�R�Aj� �BO��k�����l]`�!�p�O��+�K,�"(��|����s�͍V9���7.3���q�L?lDX���{�I?�j���q3��q�y�o-y�/:��YJP$l�H�)�8_����z�����Ao�ǐ�N^~�E�o���vYH`�k?I��U!�r�\_���ȏ&�W6���Fq�����9iV���Xt�"W�y>|m�nDpDO&x���f�_��fkZ�BM�<��_|澓�8�*w��P�=�Э[^ �
3�9+:γ5�9b����p�Ƞchk��tA�<H�Z�_Bd����	�=|vBZc?�~p�q�q��ݍV����E�&���I��30\U \�L��nFN����F
�ճN�p��$>J�W��D[�5����i	o�TE�]�MͿ�����D�}}��D.8�����!�Ҫ��� =((ܸ�o!|�lZ���1fYҘ����yY��b�΄�!�4��괱��

2�"^~qe�f��myE@�����2i����ݷ7�ę�It	/v�0�#R M� ��"��n_F9&ZZ�}�����\rKB�V{b;�Y�d�N��^�������6��M�V��:%؄_��bo��Bz�v؇��Ґ9�5��u؊>2S�Ȗc�E)��F�$�K�&��\&��#��e��	!�~���5!o�H�i~�.�1����$܌?�,�d��r��q6C��!��L��*�<���1��VSE�e��p?�Uf.���U�a�f;ٻ1�ɰ�h�`�� ��a���Ü�=�����`+b�C�
�uw�]��^c��`��L������zJ�BpbɊ�v�^3zL@[)f���Q��G}עN���键F�����I:�Ǜ�أ� L�Q�1řl��i��~-�w:s��e��~�(�9/�nA��Ir��N��;�%����+Qhq;X���H<�B,w�`��2����`0b�#�t]<e�+���]�w&�\M��	�r��Я�Ђ�ʶ�9��$�b�$�L�G������'l��dOˈȼ	�:����v�ڲjg�z��D�ɆK����U��c�s��7Kk{�C� ΌԭC�ԭ��~j���v�򵘴n;hc�,i�ik�ۨʚ�V�En�*���_o��%���=�X�(�k����F��
+�d�J��\ں+�\�Ԩ���e���|;�1�u$��]�_�Dxyv�zD���Ᏹ1+�Jn^���M�/S�������f��'(��:���-Z[�+�K��ҖA�\C�5f��q.[HQ�{	=V=����}�����b���T{( 4���a�p+�E`߿:�_�v.�ٜ<iά[���m���4�?��F�RZO�hl���pFT��miS-X��� �?��sl�7��'tJ�u����Z�;4�uyW2.�	�F(�9j��"<x^*|R�P��O��$c��n�_��� �p� ������I[Y�O'>u��ـD�꼲Xj�}ck���5��+���X�^�]���ئ�pP�:���v��n�'H�qT*γ��UB�h���Ӗ(^@�":�y��F{��hR�좂᭾��rJJ����&CrV9���=���+T�}n�&��E�$\*$�g�P�\��:�`��0�W��U�>->e�\�?�b��f�����@�n��n�Å�Ce���u�o��\�����l��-�wk�tk���0t�~�X��:{�]��ľ�}�5A(�_���B�w���{�D��޵�?�q�h�U,v���a�e��h�a�sO�wK�$ WN��zrcB�`���sN���{��P��h8�;�j�WtˏZ�Բ@��}9܃X�� �=g�OvoP4����,��
6��J`�]+�+`��n	>�����>ؿ�W�*�"t�F�q����c�\�&�M�/�d�n����CM�t�2z�9��aL�D�ʭLD�$tj z1�H�lpj��:8 %������ju�_6��=`�!��hk?}�pp�\X�c�2�`�N�%_ -������03%�*�ٮ�k��H�(�dB�P�P��K_�D���Z-�k֯�Q� �.i2(�ezaF��/�SÑ��S)�Ɋ��g�0�Y����ڵm����a�;�hH�{��\���b���#g�6��L*�dU��X�2�F��?(]e@θ0v���0tDK���߯mJ:�(���꼣1����d"~�?DN��4I���|#��z[݃�OZ�[ +!����3���S�T%�N��H�C6s���]jm~�M�mp��� ���9�n�ޖ���M����z�~$(RC�l�0u��"$5��}[5�s�?��-P�ɸ�����(�qe���t��մ�0|h��F�z�N�.ă�J,�ӱ��͋xp�9�(��6�`)����Z�.r�����L�5�q���g%�݆Oa���Hq������ �8��}<��0��OY�R�d��C��ĹǪ��l��������A�!�����C�P���xD9�m?$��_T�@��Q�¸U������G����Myy_����u8���I�`�Q=����}~OF���D@6U<9����LEf����.��(�)���`���Ky"d�n� Ã�����\ݙ�{K���M�hB���KU2�<K)�������G�8���r�'��)$~AK��q{b����A���[��>W��b}d�"����a�Q�v�]��t��s�#��F.��W�ܜ�q�D��l�s}(��b"J֑G�Ia�,т+���D&������CxR�c�)�R9ܧN]�C�W�q��&|2*Qz�H�FG&R�m�)�4���m��My�5��Ը�n�ƈ*�H�6��t��R�?#�*1F�9���!U��:fP��/��X�kS �R/���t��#�y��z@' Rt�=k�3[T�)N���1&�_��߼;��.����
��~���b)[Or�!����r��C��2��Bc����7�P\�E�٧W*�|�n���D �xĜv����8B �ӡ�r�>���*U����C~R&|hL;�_��v@�@�#(y�>)�P�ޏ_\��G���e��b>�By�UOS~I��Ԫ��f���(U�T���r²k�V�dUń���ȱ]�v8�E𗵚P�~} �� 0F"3,:ρ�I����l��b���9�B����1Z�׃f|D���Q;i]��
��oso�^�{:�5�����66�>�cG'�K���[)@�G�1H�K	�4Ή┹��>���^Z�d*C^H���P�PT7Ww?����<��H�U�Ch���y����ٟi��������b墌�A�sQ�V��EB�����8�S19K����R`�|_i��/��Q�K�Ӧʨ��� �ҭJ�ݟn�8�Lb��@��E���Km�[�G��g�@����@�%��6��8[�FnV��
F�����N��<!x�:��#J�.�=V�5��Y��C�{*�n�t9�I*k.�l�� !�_4>��p,NT_�A� 7��@U;2�xy,��W�վq,Uu�R����B�����2AvX'{+�3�\���P���qc�^Nqlujm�ڡfи���Po���l�`eC��4%�	}n#�^��`�T��A��ݧ{��.�4�4G# �ĘZ���P��T?W jc&I�{�����lJy��H�
>Z��o^`Q�_r�V,6�/�e6~c/j�vDC�`h�@ڻ"�Za���`�:Ru!^$G���%XuG��E<f��:ۥ�8g�{rf�2Y��Au(%�������<:ȉ�欣T���Ѯ��r4�$w���{XR�5#D���%H�(�E��΀��Ce���f��j0,��9��k��?�n��Ym��'~���ĉ4�j�[�\Eq�����mj�����Cԭ���/�u����FՖ�5��� ���o,��in��o��i	��T����������2��#ӽ
֚��<�(�Q����'Ax��Gd��ܞ'�"���t�1"
���6�+�[�%?�!����h�O	|u�.�B�+Y
�`�B����T��̡��(N��^t��݌G���= �1!��TfV�,_cG�v��'A��d��ڣ(C�3��fF3B���>�,�&�nv�(v$���[9����B��Kq=c�f_eTN���4�0�Ht�SM�9�40w]��>o�Y��
��o��H{*�5ʸ�U+�O��X�f��s�֣uٖQ'��`sT3����<l�O�"�+�Z�x�K�н�vN���ؘ� }
����+)�:��m�����C��kTD�p��c����͉Ӗp����V�➈>��;�<��3���@���GW�95�<^l���I�T��UcB�-Ž'w�.x:I�S�3��F�HжH�8F�b,5���]�eo��袅������;(@�O�������!j������׋_��cK�����$�vd��-\!�u�c��t����a�;��+�(�2��f�˶��{��H����"z��;%R� a4�"�����p�ċ�Fc�o�,�q����j�����Q,&�!s��WR�M�:u���
�u�n�'��p��j뉛�3J7�N?Vn�;���y�ݕ=�P�P�J���x��Z��0�T�I�Ʒ�� P���Ca�$��[�b���r�t���ȅ���16S��hD�wOOM�h̂���Mhc�!�� �9���I�6���m
���`Q��-�&����d)9�gu/L__��D����Q:��CH�޻lqG�)n&k��+�4�����0�Y�Y�	��h$�5O�PW�I��H~O�"��,@dH���^B�m=��zߺ�`��['O���M[z��b'Z����|Q��ؠ>J���P���n��P���)�!��)�=�J��yrV��T5��Gma�U���썯�=��J:�c���[wO�E��	i�9�w��a.O���yr��;y���Xh]1�^��^��P�p��XRv�ߐ���}��Ф9,�%i���Dq�<���E�7G�π����#�R�.�:CQX�O� �k8N���bG<�BkD���!���O�	�5�呬 �3����C,�DHt�cu�3��(�/��G~v�H��7j.Z�+� �.�*s���)�{�� �	�E�Y�3�(����<�	��^�\�_��Q�F��y���B\�
,Ε�Ȭ�#Sh�ϕ��b%�N^��B�Q�RX��-lD3��R�k@�	Z�͠���c��s������(+� O��/�Z��C&!*^�$]�efm�H����c�Q���H5'��c:���DU�b8,i��0��ۭ$J�Ɓ���l���m��U�����\G��^��_�V��^N��i���-�M�S�v��_ާڦO���nݰT�%ʈ����j�b+��`y\ ^��f���P�
�s�eẆ�	yEN���P(���}Z�"��#�zi��Q̀q�y��KA��.fNf�&�у�L�Bm##s�n��6�.-/ʪ��`�-��!�<�(mvG[��ֈ�߿�OZۨZ<�v�Œ@-�b�����:C@54҃���D�Dж<d��:[ֵ&j]�WE`c��	��y��N��MO�~E�9FL���"��GtV���\�ڧ��z^��o�}�m9�nGq��5��B��n%ex�WH��=Պ�zr��O�I�S�A7������Os/P� 3.\�����Q�fDc� ؓׯr�m\�׽_��G�9*g#��sG�\�-����0�Ʈ����1t�<>2rC��{	/ST*4K�<���w>��T3�h�B�B���`���ge(�$�D��0�GlRxl2���Jg�"�h��1��B��!p/�S?�N'ffs!�fA�w�w�\��;�/@�C����wW�Y�
E��B����&J|�]U=��E�b,����#o_}Ͳ�R3Y�kZ��ES?�[έ���ȏx@#��/o�Fmr��[ਕ�+���
�*�"\��Њ�^,g�_�/n�ė`r�bH�z�'4۫�7�b�{��)���̃�us��!�d��=H΂���ۏ^�9�'��z��S��&�r��]ؼ_�,�}�'?�)̋�]hr�_d��)�������,\&�|>#h�L̴�eų������7�9Z�*N�(�_����^X�-U ?,��@8[��Ş���Aa�]lP�ZB��u\`�p��9�T�E�Ɯ$�`j�yz̶�y01F��i�,Gp��O�T����à�-�K�
lϴ�"�C���W_�]���6DpB���3f�H�C���c
��FH-s	�?3d��x1���U�,4T�D�d��*�oc�G��q�h�oS�ˁ�9�e�vШY��8�u >v"yG�dE�}�zN�2��4���#�����H�h�;é�A%�"��=Not�ҥ3ٷ]1�V���"�e*��;��F.@��{����-�*���O1�d��n�����X��;vб�M��?i�Xx��w��'�ݔ_�!ʔ�lh�hoKVɂ���Z1<�e����p�tV~J��}�O�ƅ�,�Kh��PB�s�k� TY;���%m�f�Cr���j���;?�`}�K�b'�sy��
rZ}�u��z�| ".-[�Pfo�⃘`��"�>bB�-�a���L,�@�܂�E֚X^�K�f�B���ۡ�mO�Z����PN��pIA.>+r�k�$0�Q�Έ�>��VtDȤK������@R]��������πϖ��-��ڵb���e��fY�$ن�p�����v��D��è�k!��3݂oP�%��̑ ��#�����=W}�Fl�p~k�W�1J��������W�%j0��=��X�7�swr�:�*Yo������G�7������ܫ�v��:	"��1y� �mt��r���,��&�qt<��\��TN� �����$�R�iXy��$#3��0�G��ao�k�nU�C��"r1�'��=I5��	 ���8�r�E�p��4��l,ô{I�n���,� =�糖L�-bT`��s��;w�e�m���r4ڜ�'�Dic�9����Zƭ������,r+��z�c��MS�"�aw"i_�����I��:_2(b�"T�cY���YJ���K��U6��ɍ��L$�-(�kOMg�1�y��a�zl���
ט�l�˱�:���}��]���EN���%�1���ʮ���2p��E��z�ބ!�}7�QFbo�8#�,( ?$,^�IO��7�QQ",Ҽp�	�y�>V���9�U����I!L��nXGbG����V��l-�jE0U1}�4��zzǦny�[��ߧR�q�O
��A�+H�L�V�S��Z�V�`�\0�F�Jk��t�k����8Y����YP��H	CO�~㘝]FB��%jƲl^��9e�
��ܗ�^�p�Ʌ-#�F9)e�/`�:y�wiL��2��0�&|�?O�(���.fA,I���I���1#�#�57�VJ���	�v'8�w)���syF����m������/�;���#�x?��m��"�7e�b��	�l�O��.$�R�8l�Y�յ߫z}t/D[����F�=��w�/s���^��"�t`&ס��K�{���Q|x��-6�`04�˓D��ܫ\d��ȭ$��W�P?��/%��Q��X�c�D��1�g�Wp�u3�J��:���m�X%�8���r��{�"&��;��RP�s�TT������&2A/w���<@E�55�m:��h�y�z�O/�엵 ]a{|M*�/�N�cFWM;��F�g(��bA��Qk��({�-�F���f��"[��4Y��ˇ~b3�Q��=���6��Y ���|SH��ؽ�%�f��n���ð�_3$ݒ�5�\�L;&����v�S=�f�K��F���q��@'���r=f6�_�QL�����������w�)�}��)���)3���`NC!��j�e�p�hu�F����^ҳ�T�{���IP"`"���Hӳ���c�AV�)f(%	�j����/�As�(���ǯ�3��nK�r� �\ܙ��j�:>����l�IHg8"�����=��LS�F?Q����1s��4rן�P}DۘE�r��@.P���ᨘ-���.A�I�x�i�R��Y�B7"!?xΏ�/2��⫈�I3�C���TW�~B�3ؘ*����DA�/��\&L�����T�p�F��g|�q&$�w��;[�ԭB3��7[6Db�E��chݯSj������7�*ڒ�(��o�)��/Awr���3N���}�݆��0�����Ō��옽��]/IEKn�f3�E7�������n��z��+�Oہ�:+&9+q.�X��D)�N��d����<~!"�����Ԣ�jϢy����zT���o���7��4{��N�-)���T޸��D�ZxyY\��eQ�;7P�� �[\o���1ŧ=聤_�6�w=0����H$�#w#@�Z�+m��<�F�P�i�f��lʣ��f��� �o���sa�s�m�)��󿐵5�;-f'3��w7�����T+5�_ةiʻ|%;�`�n�B8ه*�W���@S5�c�\��}X�C�Ô¦/FYa���|#П�L8��Ꜻ����&ݠ��<��M=ظu�$ͪ�S~��g��b2�?ş���0=�r��%nؑ�?-__��x���(K���K��ރ�>����,?���yF�e�g������aе�b3h��Kz��i!��t�����/��Ii.�I�)O�+e�^�\7�1�NН��M��NS$�e���n�x%ꚱjb���нg�v�`��Ц^H�@:aa�=yp[rt@B�����|2"���������¦�f������_��S~iz�t�^��*t;�K�B��?:���e.�k�JY����|��)!�X'z�Fڕ�A�]]��$lfD�{��{QE���_#`킵
v�|�=�*��W��f�;"JN����ug���2g3��]���8�]��嗢�J){���@�~%��s�:��0��mw��Aj<�� ���Bu�W������}����tEQխ��>B@FaS) P����_$߸��wY ]kw_宂c�o������@y���	�Z�f�t�B�6�" 0N�)��S�gk�����48]x���dS�����gٟȫs���bn6�ǣw�02�"_ػg�;҇�VJi!�6��=X
���/Zز��^�%���,��w2� �I�QHB��ZN�Sk\�o��zE�f�P)Uܑ�e{y��-ؓ�g��=�;�͝�p���楗���~PY�q@�w���m�t#����,(���׀��o.0�y7�8����S8h�>����>#�q�?Ҧ�� ����%
�2$�ә+ab})r��%(J������2T������(1���et�z�(��q̏�Rm�(36��P}c/��P���Ӡ�u1_�r��:�CM�e.�?p^�{J��|YY�	sК�Z1��!b~���L5{1o��H�X�	W����%�:S����~�`�;=%�Z1\hP���P��C�d�5t2R��lұ\+�H�rkZף�����5��7�I���p�]�%j��c�\�\���
]�}	��|1����.?��{�S���rCb1�(g=FW{��A��Cf��lF��W�Ixzl	��B�Fd[��H�#�j�P�n�N���5<���p�Vm�Bz5�fTx4���)RR0=�tT�<<�#���7Q�y71͇����bWD!���Ŧ�Q6������8�����Y��i����_#m�̏΍	w�T����)EH���"#�7��1�����#��=���rK2�TwT�M0��K'����h �{(J�a���ԧu�L�� b�e.Xbp�����a
c�������54�E�j~�o�-�S5���q�w�Eg�i�sG�WX�~���g�8�J���<FNMS*|cL^-���U���ГX���
�pvFH���,�M���I©o�xLYQkn�w�)4 xd®��62�ұ͹HU|��Ue��H�9l0�����$�t�������&�^��[2���o�<0���M����^V�g-ΊǛr��8іň�k��zej9�CZupY�� 7�� ��y�3w9m2�ȷE��E���q�>��.e��Je����!�U��8d?B�l�T=�PNs��[o��CL�&哉����<�˱?�#AFW�=%+�t��_�DT���ǒ/�������ً�m�U0��&���{,IA��e� PQ��6ZR�S�zF�xE;��>	���V��Z�,�I�#$�ڻB�D��r�&"���^��9�^��L�%���9^�`@z�_6b��b�L�`�^�̚c�(��Й��	�s�#���`�t�,�2x�/�!�J��Χb�L��UVto�����l<b�&@Ӽ�/%p�$��v�� ���f�6iI���^���s�N�m_��Ɣ�_Ս�1t�����2�Q�fCr����̗����[x� �;��1�aB@{�V�2��[>�5��K���4���&I�۶����[�(�	�eؠ[��<��I�Wo�y�pF}�\H�,�;��'�*�K/�Z�����b)b3�ԕ���ݲZ��ۥ
�a��aD��yЇ� ���mS���鱚}���ԵJ�}n,�'ᬨ�j����]��*�g�=FeA#x�^>�s����н%�1鰳�>8g͙�V�uþ��Dq9C��)Mlw̓���97�I��?$�ƫ�TJ���p�<�8�^IL��-@.n��]����}C1/,+�n�K����U�6/�V�&q2����vlVF��Uc���(彇宱���}���>\����[pC:fDF$ߍ��ZX���3|���Z?&��D�Y'>2��R�R �bS̋`1������i�O�[�~t�
��X���$�4�nRdd�zu�����R�#i�@|��v�yQ�Ց���' �H19���瑆��M�R��1������"�\ߌ���0
U�jv�2:�X� �֋N�VUк���B)��L�4�
v?����sɁ��� i���-���q����L�Y��{<W-�� RM-�������l$��cl(�`�?5��F��ʍ�~ j2��-g>xLG�b� �"E��(�C�?������Ӎ�i ��X5���CLn����0r����`b�#�R��`r�帿���$�V�ꁪ{��_Jn��5�D�A5}V��t_�53��R����[���/�:~���kA�����}
t�~�ήFviq=��,�D%�zŶ�˲i��0� ��Io�j��R[2�7$�񇿳�tW�y��7���i�g���R�8�G`��j���Q�d�
e�����Yĕ�_��A~����r!�R�{L����kD(N����c��R|O�vvxa����f�#>W����u�9[�����݄�|9>87B�oRr����"nl�O�&"K����9:��th6�]��P�|;�s�=�����.cW��>$��ڡK�(@���Ѫ\?����E�H�"b;R�yv˹$����xC�i m�=z9�V2q^����KM��t�j��E��	*���0Z����k�3��o�9��B�yL�b�����Su
�,�~\����aL9��:�n� ��C�v����{,(WX�����e��P#��@̎4��fb���~�����<�G��dLJ�pz�9�F,'��f*iuE��HҼ����d��D�Eh�tJkM&�*����>�'P'�M�%�ܘ�+#2.dЀ�����ѭ^mpѳg�\kW��<JNT��!�bM��72_|����WO��'�?����Y! ��&�_6�� ^����6��cKr�s�f��W)�J���1/���f|����`0�FO��cC�"~���.�u={R���yde�4(R�����	2�7���c�)p�=���x�q��(jk�[A�7>��Lrb��&�=C�ar-�g����u,����C7AL1����_XVqI���>����<7����q�����r$"�|�i�LS�;���:���{��zK�62v{��Ȅ�|2����"L�O�fϪԩ�ϔw;E���M�S�>	|���3��VU�6�-�um�ЊrM��_���ݬ4ף��?��n�U�E���a!��#���?��Ý�?^k��u�V���$�n������̻\�5���F���耣�0+���x�U��|h�ǎ�jC(�5~`���@Q�
9���i��a�\�́��p�jJV��\��s^�_L���7��SU$%Y�O���st��ʿ���k@&�� ���<�n�&Űߵk��h]�	�pM�X�+XQҏ�x#a�eӸJ�1�9p�}�r�#�Ύ���B�?��*Ja���@�S3��T�jL6`Xx]�JVQ7�q��{�=S3O��P�QT�l��Zx,_ߵ8��ʒ�}� z-��iL�24����ղ��W�[��`�4�e���}Fyr7sS:+k�������� �F��h��̉�aЌ���������Ƥa��}t���3ĘR~���;ME6;�j�N��d�9�����d%ۤ���7��6�Q�]���&++2���U!�!_�ʬ]��*�Ue��ظ���o���E�W>��Z�^�t"P�1c�i׻���r�p]�LP>$��2����:)�r�,��^����ak��6�������V$%k���(��c�����H����Yz�U�^!8��Z|����H�j�;�����1���D���P��*��[�;�np���ɮ7��
�WH¬&S�j��:
W��4+�,ܙ��Erҍx��:"s`o��!�`��h~a�8<��˴�;�O�|H�TҼ��fj"�ٖ�(|M"m�{h=�Tύ/ڞ�j�,	p���4�rVxmn��!
Ú�<À:3<olU����F}���_'�cW� �Ud�v�e��f�IG��l�#4��h:���!��w(��g��[�� ��^�PGv�R�]���F�_�{L� wq2	rp�v�'sRc����R�:�jǛЛ�������:Zn"����<)+��*��i���~�T3��e��e�c���'jh��Z��S��<���s���|T����8����rq�l�� -��u�|g!�����T�Mb�_�u���on!��jxp"�:Z�Yv��o�Gg�������;��^ַ�����P`�;z{��m���NV<U���Nay�.�̚�T�6�����?����Y����#�o*7^.�A\����NE[ #\)���Ō�)R'cfhS�����{��/1 �`d�x�`��Ey�~i��KƆA�.���I�^K��L�3}�JPؚ�q�fq�g��a�w]��ؗ�. �6�׭j�0�Sʧ=�ALMAse�4�8�̯I�ƃa�5A�y:*���,��z,��9�J�ɔ�@&��w[U�6�̈́��n6gM�k��A���J�m,Q	�*:���sj��^�0
f:�]@��^4�\����8OM*�br�)��Ѭ�cZ�q�k�B�a݌|GR���.�w7 �ׁ�6�Q��Hf���+[Z�'�ZQ�1LS�����4X���^�_��*����6l$�'C��g�����f�=j�С|m۰�,��,J��<�o�WP�5;�'�7VM<q��g�ʛ�)�sUFEc��kB�M$Sy��t�xQ&�W�H�z�e�zFd�`Pa|�n.����ܤ��k���_"&�X룆�lR���j�)���BJ,FY����']r�g��5�fNl��0���K���N������0�c�2W.G�MmV�V�j�hk*�N���ZGQ��f�~|�a bƑ�|9J�Y1�{75W�/rZ�x�l- 4�}�TC���9�>��	V�+�>�+6�J0>���+f�4�B��Q���j�"`32m��-�G��P_���.���@/�<X�&q�{�����6��w�CQ�5�\�*M�?�#pTġ��ܶ옕��7}�;�V� R6l�����	5����OKJ�OX({��f�}����c�!�o���ښ�1�D
����U��	5	I�dm�	�d��x�P�[���`Y���X��Y���٭٤9/�n�(X��Ϧ�G#	�Vo_��t&�eI:j�f�K�G�Tt��k��%�Υ�
���n��O �����Ϥ�@@��w��/Pa�(��`l�өZ@�f5�#U���9�r�OH��Ԃ��$��`�?k��jd��CCY���"��[�N �˶V��h3���[{�Z�5q��1IR�9{	X�:�Ґ_�k^ʾrW�W� �h\��
�d$MшųV"U�i�&!�<��͏x�oe��Q�Ո�_�i]f#��ی��OP�I�2��b�H�D}j�K��&r4�N�?!��E��!�[�3���'��k�3ӫ��	���F��6�l�����N��U��3Gb� �51�u�+agTH�L�����	(e�0:��8`�v�S�:�5��E��1:��Nl��#��Q�F\]��vM��<��9����j�R�gai�	��֤�x���&�ȫ�{�?r��i���Q挙��D��6�(� ��9���Ic�h
�>/�'srS�R]��:[V���s	��>�%��4 ��Ǔ|� 7�ێ���4B �\w�A� uAQ�7mx�׹��s�eE4�_@ {�����Q��%���.��cU�_���s����@D_h�,�R£����0�ݓ�v��p$#��$T�N�r+��ˊG33�k7u/�t��}Cc�OE����"RC��<��R)�5kl��Ys�Cz��l4����������'ް�7g��K\�5_d� 1�r�9�ӈb"eJ/�7cja]��ɡ?�\S�^z9A��d��p�1�B���uyb0�]�l�^�����Qdf�?��M�dEv�s�[��%IYia"9'�¶FvV�h��"wpHc�,�,����V�n%}�pd��k�yD��}� ��*��G�YɄE���4WuE�#�e.�_�'�����GP<:�
�h��F��[��x�7������nW��u�C<g�å�a�5T7N4㗬x�N�~�xk���}x@�E@�I�����fv�E��Z䙻[�a�<_��ooQgL��C%͍�W�q2D��ŋLGiK�e�E��;
��-���䝶�:"Fb&^�ʅ!-��P��{Ӭu�MD�����^Jb_�[�����o'  ��3)���Kh��(Ծ@�sD�D`�����a�'��1�qQ[\/����aoH^+�o����a���o4��Y}��G�����W���Sz�j'n�
l�\L{���"��\��a��M%��G�%�U��aR�נ�n�4��]���X1�?U���c����v�Jp�P?�f~��Ud�63�u5�h������[,O��,$��&Q3��Y|E�w(�=��8gJ;�Rۥ���J�W<��A���J�iX-��E$9J=
S��_��MIp�ۥq�9#Wӽ�P���I���II��^�Ņ��f���`�C")�/Ω�7{-2��U�������#�z�ћ�ђ�L��%3�����r��0��\�{^��#.� �<��q�?�n��y�@M��y����,�.7%&�$�O��e�'�>.v{yU/���j�"�gY�����*c�NH,���^�(���`��u�m���
2����ڇsv�c���Hh��0Iv�$�*��Y1�;<�o�`����v&�\vԿ�Č �T�w�E&l��*M-��y�5_��Aż��|��r�KQw!U�%y4��QȣW���I-�g�cVR���|z{:�ْ-
��1���27�"��je?�m��n@t��m?s��h8�.ߛz�ܣV2�����������)��,�o��9o�x��h49La)
&�L��g�� t��XZ�t(�����_��+�-�m=����Co��w1U����xNҿ�p�{�t�5�;&��{�nY���s�Lיm���5���(�S��6Y]�d���.��7��zn�jG.2~{@���(�&{L����֖v���vm�QC暙���&쁓/����]Ěj����#RU�:��م�h�`̢��h�s��=�N
����4ٸЌ�Ϯ}�g��]|!�q"~ӷ�*5�;I6��`����^�����(]S�c�M�V{�h��sB�X�Q-dMX`�p�M8X�)�S��ouCj᨟�Nr��W],���S�ܪ@��n������ܨ��ca�!����O��_jIܮ���({�z|{85h=V�[�@����MK�^���"��� �w?=x�c���mA��s�=F�� ��P�I�Wr�����Qw�e� ��PhV��hO�G�|���Ӈr$��m*���H:���"���	0E�s�j0���������~�2oi��˹�njo�uk��N+����S0c@m����2�Őڊ�An;}�F�^��,�N���3�䔕d9�n��d��t(��@�����{�&�k�K
������iKP���(�G�|��Q#�������!��>�\"����8�n�,%:ie](%��љ�澼��t*��^Q(�L}��l(�چ���Q�
�|tVB�Ƨ��u�H��[��`������gH>�q"�]Ö��'��� �0��K]��Y5ϳl�(�0w�6XJL�n�QCy+q��!�W�ёE������0T쀶JKs�tP�t�wΗ [3t�7�q7�<�/�?ۘ��wJѕ9��o��de�R��J�L"��uiT�w�x�k:���F����g���Ke�[ ی�����F	�w� mc��tM�g�M*vט�)'���;EX3q�6{ʂ/�f8�fYȴ���֯ߨK7{i�y[���D�-�\��T��CF�����?��Z�n>ǆO�t\�;S����l�T���Ş.�lJ��by��X���1�+�
mO��U��3:q��������_���;�r�V<�V9G��B��<3v?�ΥoX
�&�����F�H��
���v����:T�O������K�#�9S"O����iFʕ�	.�4�zb
9�Ӎ�,��.qO�K�|�+QG	a�ੳQXt�jJ���|�s�h��_!R�f#��gXq���}��vK|ʾꃈU���-B%R"Q]o�Z�S�؈}��u8�]�T�z��sm�K�,pr��r�+y܉����;�3΂�'%������$�聞��$�\  ��ǂ�g�P_�z�R�5�oG��Q�a���\�`M����n�㬸6��o�݈���hTC��T[���8�Z��{�th1t��q��5��].�e�]��y�U\�������K�鷈A[��0�H]��t��������1�S�l�PR��5:x�*uP
:���0#�W��'��&f�Ov=�1
���'dJ�2��7��W������.�����;B퇣;��\�"���e>��W��B��c�Z�\�/�c���K��e���F�+��	X=V 3nw>Bre���Q�Vr}��N��	�f7|�������]��$�C���8XN�8Ƶ�"M9X� �-��V&��F�/y�C\D�7����
�t�2�)���&Y6z��O�����
�z�2p�:�c�4NJ�k\����X&�"��fo�=�y��" ��!��	��NN��+�6�]lZ{���ıP�����ɽ��.kx�0�H�7p����'=�{���@�Q�f���g7)j��^2�^3o����x�.�)Y�^ B�p��ꤗ u���#���1'цRȣUѲ"�]7�C���Uo0��&QM�amjk��]���8�f�za��`=˝�[Ծ�pX���-oP�^�d� �J�Pq��X_���qBA��'i��Z|R"(�����]X�_y��K���㘉��M��G��' `T$�� ��� ���0��I�f�����<!���<�ߖ��::n C�r����~���*�;S�3'��ԉ9Uy<�p&���/Xf�	�>'�rt:��#�*�G���5�É��c݁0�%�X��?R
�R�����Wd,;����Q�mFd�V�E��;�2b������~�cи5�������LUS΄>��Ԧ���0�+b��s��Ř|���{�3��5@��`�Yb:3�gi�6 ��.?��£'��_�7Jx7AK>3�\DbkLI���:bk���9�.���.ʑ����]�6`N�z*�Z�Ү�����5�k���u��)���B�m.6'@iɸ��͸�"��wAⶡ��W���!�����V�W'm�R���D��@��wj��Js�zgR�c�8"䖏�;n}Z)~��i%D��n���b�c$��po�-R��{�<�%7�P�ʲ�2�ެL�m������rK�#�9T)'`}|ǟ�?���`����G���넗 �����m����.�u�y57����X\��w��x�c߷�=k6 �r\ �CZ�W����A��N�y,a�ޘ6�m7:k�~x���<�:��#x`Kb���V,.R��G￶����(��{n�,7�e���`|�֖|`,��$ B��w��({�
w+G��pO���r'�h�7�*)6�5���<J��%ё����c"���?ɟO���6&X�/����l����՝9�a�-��p��V8*��E�V�=�gs۞^��t�2X#�Jk��UsTu�[T2b��w�^.��b��L���t}8I��{F�t��zź:t�0��r/���z�m�(B��rP��g�����l�s����'癟M-�L�ʖ��cb:��|��5H7�ʹ�E��]�#h�:>��ϝ��ct�k�^@f�7�����7�J�o@�5J�|O�.�~&A:��`My�:�Cl�c�;����3����dbbܹ�۩`eQ�ʾ%wݡ�Iax*6���\Zw��3L!z݀>z?)z!ҹ�@X&��Z2��5��������{��O�)�n�*�W�2�Ī9�e���d�?��B�/&�=P��X������k�r���8�3hG��d��:������L&�\H��c�@7� ��AѲ�����%�՘-/(���#F�C˺*����O*uxq�tt0��6�,��c��X����Q���JeV�o�LM.�BC�������Z��h�2��yᰶ���oħ�W`0��#���<謏��g���w�8,H�P-��C���@���EK�M�y�n&E?��r�%��u"�}u��ҹ_�\~��r[��'��?�c����Xk�]A�y�Vi����!�19��y"&ҘV�[C��nT[�h���9sf"F���{2j�>��|\Lul4x*�Dݚ]Fѳ%:���FRJ����\p>Q��K��&�e*�ƜE_�h �	�˘�c���GHЩ�0y���?}��=�6�n�~��qm��vt�[p���VN{�i�_��u+��*�vq�/�Q(��hU	%��S?�U�0&M(����?RJG������Dc��v�M���9�Y��ydG���Y��q�*��I�j�<�������'�4�-fz�u7�/О=��q;����S���`�/���<-���
�D�� e�N�c��LF��SXHƊ!����
���Ψ�wZ�|6�g�6i�Z�|���1Yi�*����o�慄4db�p��(AY:�p��V�(5��h��@������q�2��*J�B�?�$�ek1G�dZ���/(Xy{���I-�c���Ȁ1�hi���F��<z�ݔd9�'P�+�͞��7���K&c�@j��~�e�7�#}k�$;����b[փJ5���)�8B�}
� TB{|��YD㐘k�c(���V�̺�����Of&�Ͼ��bT3���Ð_$}���Bw���g�$�ifL�aP?<�V����g�M�v���/�+�	�z Vx����<\z�.�y\�s/k�iz���"*j,�[�a	o���sz��߽�[�v�Tc$ү��\�d���3X�n��}���#�����0D�D�m} I� Eü�0��\=����k����*�6Ƈٰ���޾�hw�v?���h�A�B��A����&��EKQ���d����wQ�G�Fh��)I�֜�_lZ�ԍo\����Ԏ�fz��:f\|�����%`v0����t%8�E߁��+P�3�'O_}Y�����[�l�r�i�ԝ��c_�\^ �w������̷�^+����u�J��������&ɋ�gQ
{hC-���K�ZߡnՅ��jw��D"���iW���l��Y�3'�"�A�8�ɓ��}	�GB�۟�ӱ%���0�[E��P��=�@��W��d�s��?����_��Di.hH��Vfm�D��u8�خ-ŜΘ�Зq�����R	Ky��f�~绘V�H�����E��Ikn�6�b m�z�*��Ͼ���X��ђ�d�������]y��cV�5�{ד��{ �!~�K48n��:PJ k}P�f:�NnPY�xW[�,j<#2��<�hb��8�˨�x�B�~��+ε���h�|f���,9vn�� �X�7P!Bf��w�_�+��[��U0\�ڝ5�ޔ����7_��828���xݺ�����&u�	�zW�GHD�y�F�3� ��������QWz�E���	Іq�<��C��*G�D��5q���?��:�ҒՀ>��dw`�3۝���"!xY�Vw�����1
����l�xnx��M3�5��R��)��+L*	�qr�4��˴�Щ��٧E*���՚��=Y8݊���&x�J����5y6$U�j�e��bJ�ns�W��Es�[f3�X�T��P��	� !E���tϛ��a�W
9%���F�ϵ�YnL��]��x�F�O��V6e�-�3H�I�	����3
|�Q��~m,���
?����!������V���d�(`u��o�ϊRzs+��O�Y��Zx����7.�1O�<it�����:�2��H��6��������Zf�%��dy�;'��ޯKCA��Y��Zn���\��H�k��r�SA+t�z@�RB9pt��7�9���0�ۻ8
`yy�}����^_�b�J��D�<�!~[��%�W��P�Í�����^3!,2kWn�m��A�i��.��	ҏM�i��(K7�h�E�l"�V~v�&����C�h'\��Ϛ��W�y���|e1m�"�iݢI���UNju� S�pg��!vt�V�`�Θ����fƢp�K�/�4@ttAʳNa�}>�ǹAj��!/�޿Z"Շ���52�dr�5V,+g��b�d*Q[�av��z�\zp�YjΫ��.���#KL����5�
Ѩ �����B��(F=��m2ry�7�d�R��a���$��*�)��ȿW��D*}/�H&G�>�gڍ%�y	�&.�Ņ��G����]峹�{�Ň�
�����tX+HX���w̄SxŚt_�"K�����z�|Ƶ�Oj�\^?h4"��8��I��Z�PT���˝g����S���;�R�O�@r�,���v��r5��b�2�-3��(��1�$8\t������5��s��=y&�F.�住��������/,j���X�!�����Fy���� M��"p/��&l���"��n�R����P-rgS��	A�L` W)��<H��lHȗ��#yA2*��L��%W]�N�I𪘫�)a2�3k���r}3�6(�&JF$q	q���~I�F�d���?¶i�
����Z�+��� ��d$�I\>]׹/2��������Ǝ!�|]��e��o�N���s��s��B-@�K#�R0��I�^eXN��d���Z���E<� x�/�k��,F�_ y
w���f����}r!=!��Yɋ� �U�nO���c��t�df�+���vj��ܶhR��'��y�b�;��X��#"�?��$x�{���I����c͐���ݐ��;��e`-���>�ð5�D{��-ʑ��A�(�z�G{���35mZׯ���݋"��?��-H��b(�ӽE&�髆T�lQ�\z^�`4�K8��ȷ'�C����S���J���R@�7���~�a5�2�GY�,!��*��g�n�]���[|\��C����~S0��� ��]Wp�h3��H1�	v,��2�� ��e0~3���z��H���Ǵq
&��W�:��Є�n4�l��tA=琥/�J0g+�=a��x��:H8��CK���Zs�`uƪ_`G�^͟�Rp@74'��ܘՕ��;G�T����9��}I�[g~��wX����p��F�i�9�� �~!|�sݦH�����їT��jt)5 m=�?��;Q
?4 k�����6:,���΀-�^;jYi�vTo�!��E8�o���J>��r,�����*����6F������p���t�z�c����h�%��FQ����=5)W�m=:A���`�X�����C�6��.C��=Cwd�5������UZn��/7�3Y�����ӯpz�p�F+Fµ{1�LR���
��'����.�9���?����Aa��ib:!��HmUu���=0A֘N��D�.�r��T�_<�M� �)����>�mt��!ˎ(����"�?~����H��	�}u��-w�.;P��w��� �R��h8>�NK�ŚV��n�:�p^i�~9�W�?mZ��d��M�-K�U�§��"�P�i�v����$}v$1��>����;�`7��>��?[)�*�\Yry�F3�E�űqk���S���k����q��~I3���_�EY"s4رf�P���T?���TGE-�� �>́?𮄤���b�]���ꕖ����BY����Ιw�&quz%JA*�~���G�֋���iC	�h��ƿ�d&F���X���G����}�2�A,��6�S�E�'�oNP�ˬN����_o�������*��|����0x�bb�)|�/r�⏻�bc��	�})��Wl�oi�|��R ���ڣ�o��z+�ΗSw�
a�Zya�jL�D��*�	f��U�2U���/��g�a."eC0��HG�t�N ��$)��H5;�s���oFp$�'�Kl
�=ƙmi����k,�za��pٱ�n+�8��u���� xɈ<�rfD*�c�sm�y�y<q�d����gC>�f@$��q��W���8l�_�sz��t� yZ`���wk|'@����Kg��9��}�9�Ny���?��_�	>G9���/���iV2j�P��)B�X�N���,���q�Ey�l��S'ϠcsLqCJV���$�;�\��J��Y��.'(���[�G�e9�&�P�X[Qp��f�a�E/v�JT������5��cf�O��mMܺ��b����o��~����Dt�N�-n|$�r�$�2O;-NG>�o)��ߗ[�lV�3�cCՊC�߸��<K'1PGY�K\�;�>`�>-7�T��'nV)��:-�CZw��0v�
g�	SF�I���.M���'�ܛ��]̃�c��|�Ʋ�ٮ�fm���>�ZK_V��m��y=��Z�4��G��|�-p�f=�*x�ٶ�F�Ma�I���Ⲭl�k:T�_`} O�K�v�9\�=���3�a�r�f7��?�%NM��fL�Պ[�m[QN&=8L?��H ���#Ϟ{J��$�Ҥ�<2�3b��]E�讇�Q��ݮm���jE�r3�ŚC@��l|I@��W��^[���6_��Ė,�����`	o��0�?F���)<�R�#Y�~�s��3�c�AV9 ?Pv*]Y=����ǂ�GU�e��Х|� ����n��+Y�]�`{~Ut>0����JME��-zc��ot�hF�޹8�ʖ;5��B�Nn��;�[�7�ƕ
�޳���ٌ��`��f׶��m�W�>�ڼ��/�0���2�#��R�Y�d�0SI|iY�K��F�����A=�-���m^^�L�?F��۳YoϰY�V���!@&:�1�d*1W� ۄ��UYZ�w��╶��Q��+��ճJ窞ۂ�u�+�$����W1�K��g��q�h���Z3���| ��u.ƽ������ �n�$m�엫��șm�l�mI	��¹A&��� ����o��ġJ��
���� p�
P(s0�ϗ���8dm�����;�<�#�=6&�Pl*�A\X6ca،����T�3��jw�o{U���4V��et���Gp�+.(�T�|#�I���[>�uvBx�~>�<j0$ܝJӔ�m���O�}b��q�=`��`/`C4i�H,e�m�   �Z_1�cǚ��\�,OS�>&�b�!cq������/����l=����z��<<�")�)��مD�`1�+��7�)��@�Px$��������T���L�,�G1c�P*�P՘6�67;���F���'��)����s�c�Z�.+&9��>�$��+���L8���E���l��Iu/]����S��7�lԤ}�As�f|�K��CB��PU��h�s)O�r�&;�o\���i� �����?_g�'%i�ͻ�B�֑\$D0C�4ʶ�x�.�"��+�Z�-�S�-=3�~"�o�[(�G�C��Ԟ~nv��2�!6�Β��vWEy:�⏸��4W�z��;��4z�/"A���)i���ߜ![�0���%���>X��:#k�}�K�KUV�؊���C�����H�i��ꢞ�.R,�a'���I���Ѳ���HL^�E��������������o��~[�E����@=땠2'4J��x%9�.�s��d�ͻ�W��D�V�]��/�v���Z�п�LM���}J-]�F5�2A�4Hx�%�0��`�LS'�.
�i�H�k�ύ�����AOV�e�q�y��r��9����*!T��K��=T*���j�j�K����>�"?&���z��G�JuѰĚ��-Gvҿ��Q�Vr����	��PK^d�9�7���d�Rb��Ӳ��%��=��������8*��j
*�'����@�~DV.������{�_��ԫ	�>�2!q��N�0�FAIF]�=���W��-�Ĥ�+�B��Na8��!E�G�3#��nh���Tk�HX�c(cN�l�����!��h����A�S � �S�9�I�o�WQ�S�5�%^:J:����	Tg Zɡ>P�0���V��g�%̀��OH[5?�a��������D{o:3�v�oNk��c��(�-�~:������Bi��늀��u�(�!�e���S��+�si���0��h������Ԓ��q���D&�b:����:M�紉f4��]ʸ}����FV�Ge
�0��-r�*�C��Ir��玝�c����|&���E�A7U9�����Q�f;!e^/UI����7A�:U�Rl^z��*�!=Ln7W%
��V �,.���Ώ��'�8���{�fT�_ҋ�E��   ��	;�(է��*�6�z�?y��t�Va�(v��P�g��u�/m�R�=l�l����Կ�5��Y96�J��,XW�����Ǣ��է������)6� �Z��T47-�X&���k �|6�4�AFd�^�����[����T�d�%� �y�AR�f �͠�����$d�DI�'�_�p�b���Q`��D��,Ԅ��Z���_� QW⻨>C.n,T�ݛ��>|7�b�0�7���6�[�84w��\͊����PK|䊐��g��������^��ʮ��z]�1� i�c���!�Qj1
��\W���R���amތژx��j�U������h!�f�;��=X�h|��D�<�3�wa�� �Aq����S�n�	["����Ċq��9Ȫ�N���1]w�Z�c<��e����C>n��^i�)��Z�T����3��U�M�Jb	ʀ+"�h��$KL5/ҙ�4����!�֤��5���6��Ô�I��d���_��]�͈ �h9g?�G2q��/f�|�H+��� |�u���g	�Zy5��͔Ќ���bF��ٖI����m3��Y�\h�"P�B�����b�m�v߾��^޺}������GK�/Z9�O�����[�D�����H<�9y�9�w���X*�J�	[F�fU���_��������$�$E�H0��uG�1�蟨�!�3A/���'Þ3H#�Di����u��\��wl���c���I�+?���KQ�4h��!]>�pa�$��oROR�~*�E6�"�1�)��~��Ћ*-1����,�M��C+�t�R�~#�#�h�D�8t-\Op#�����$��̼3�����G������L�������N��W����_���e&�K�@>:p>־ȧe	�%��m龌1Cю1����*���BQ>���]�?�ܹ�B���{,r��z2�qa�Y\��>i�/rm��ɈL�J4Kp�E\@�𸭰<��4�\��N�%��	�\U9!0�e�H���~���	W�ee֖[4������2����>{��B�`?����C#��w$����K6���|hS�Ci�ͮC���X�f��̋�c6\&.p���B�S(ձmGBE��H,�6��5Cؼ0/������}43 �����E���>�U�����ɥ�����nq�0�1�|���*~[�����䟁�s�G�D`\V��O����R��5��e��InT>�	�z��a`s����K������y�v%|��4 � s_��x����<f�q����0�'��P�H�r�=e���U��if�wMތ�gln��Ecq��1�"��� I�%e����c�$�|�{t��$����p(�;NާSD��6��14*Owc����,�ϛ-��6-C��0_�k���`�P pn�x��$#�
�:z1UP�q���7ݦ���>,��%��u)U�*
���(e�4�)5�ǊO���
���˓���t}.� Rd8ӟ��)�`�؊3k1�[C����{�5;��;�9#�����b�M���r��l�ϱ���釢�7V����9� �m�~��r��������:����ʑ�C%�����?֍�F(��ɺ�hԣvHV@J@!p���	��e-�E�e�獙����<�Gf��;V?�A�Ů�`��z�j�U>�:>�]S��J&��W�M�j?t�Y��}�"I��;��ع����p+6�&�p1��9C��,��W
F���P���V���댾(�ی͚,V9�Ld���ײ|���X��|äQ�e}5XB�ᤘ���R���-�
?s^��<_�`/L�M�)~��]��I��)�����z,�sd��dP��Ta�
=�.E",63�D&�Z���
k*0��5	��CQ�x�}e�F[[i��+�e�<Ɍ�7�1���d)V@��0��x@����a���Hmۡ=4�i�8߽Y_�u|̵�	���3��͙^��!��D6�����*��~�@��#B��'���¨��0���-o�x����@򹡐������k�Ϛ�j]v1P�k���1�݊h3��5s�	�՚���I�P�S� ��9��V�Y��z�w����A��$�E��bhi]�ԲeI���g|kl�X�)%�i���ux�������p����%fK�!t�F��9������^}���h��s������1㱂��$�C&����b�b������p��0TN�5����|A�;��U�1wJ9� J�ea�&SF����Z�f})�."�hÕ��ek������������OV,�-ԫjA�~	�>��y߭cbmHQ/mǤ6� q�O!�d@k��F]�Ygk|��z��z"���{^�6��B�C�6(:^�6-܈g�f���@e���g��0���*����� ��y�ٖ'�3	���U�̸��
��2��e��uS�d�X�h�됸�����Q��Z��|���l~��Ij�@��p�w
���,+H/�Y�����L/V�2�&�g��vPX-U>�^��2Ny���0;�~�Q_ǳ�ǯB�Թ`���+��p:S�ǿ���F�>�UM�OL���ݾ����Ƿ"��'#Aam;)uJk�g�0Ld���.��tr�y~9ɶE�C�_���|����i:�}������`Z�*�c�DϢ���8�ZZ�����U�9Ӊ ����QĈh
��f��'j���+��{³u��b0?c��5�j���i܈ Qh��Ta��ǻ��:��~1� \	d��.�|^~����V�1$�}��|m����
��)��P�v�P���;���@��m⾓�w�z�Q:�-�ؘo#��ũr��x$K�ޕ}���;�*;8EM`�	��Lx���!ⰘS�{��O4�|m�Brqo�Y֮��d�iY.6���t�<�z��U��c�O��\?kz8��E�iDL���/3~ρ-���i�C���ӌ�o1���2�1��(���{�U�t�B�dv��0�����R�	�{���m~r��sh����<���}�,���敟�B��a%���Lc����R�W7F��|q6	��2a��� ���pvgVP$���&Y�:��<���V�>ȗ"��?������u{Y�[^�a?؜��'3@ �{���,�A3�*54���/�-)/�6�M��QB<��,�[�%Qw��B�7ۚ!���]���J�č��Cf�W��Á��2I�4Q�YMX��MIa�&���f�8}��rt,_��to3���,%P��A�
"�%������j�����-�ސ��"�l�Њ6<�ʃRQ�2� �@��糾*k�d?3փ����vRJ_GT��͒�+�NN�Sa�w���������F�����a)O���.�c�2��/H�?X���\�p�k�䱐���_��<�;^Ik
i�[�1�]�Џith����튃��/����,�w�ͷ�����\sR���h�B��]��
�ؙ22�q�\�Dc{9`y=�z.��To�����8֑���D��gO��2{�(0�q����n.���/1�aܽ*���.�2��"�S��Zk��k�=9o�X�EU����8���C��hD�L�A���;b���i�.�����P�ի�� }�'G�b�x��A�ݶ˳6��3M���J�V>q���ƴB���S݊��Hd�!���n���5��{���sJ��"^-��C
���BӦ������dsV�Ԁ*�7�6�`n>	�B}�
���$S&>v���1L�NC�ڠJХ�e�� :н�� �ڰ��L�m\_�;����H�SZ���?�:�h�1�0268��v'0^	*溾�
�x+"��Ov��i���w*�H�{�&Jѿ	���獻#Uv*2[�W�H3����d�g��s����e>�n s��@eH�&O�w�z�����֣�X4X#�2�CdOP?nO��uI���d���}>�5H %�J��^�Z/t�.��x�R���t��kq��~tG�?����Fj��̨� "�����b��;g�*�s�����q��b����l�aX�<���e�N�̖ws�cuJ��b�ˢ#��h}�^g��taJ,
���b��ü䰗�=��o�����#���r�o����{�/���R̞�Dne"��#D��Rõ+g!Y�{��<nz1`�(�Q�M�K//GcoHp���l�^�~�Eq�o�0�f�-u��-*��8���B��	p�A.r[��c�T��hz�}�����ܯI���2��0\�J��+]4G�p'{#�D	>hz��eo�U-J���q*��m��֝VS�q��&42"I^ppڗڬ��*{���Q!Ԟ�yQEݏ��7������iH��?��ES((�\��1�"�J)�^4�A=�$�,*iլ1��u���n�v-�+�+�+�v�����yNg��Xޕh:̸�#`�G=��aV�T�h�T����c�-��*���'���T��&�|X��5�ɶ���i��u-�*"�+
$�I��T��hYf����f�@��jkC�6��d�6E�v��vә��d�W�{���lf�,�[�.�"z�Piu�y'3G�� 
��?<�i��q�8��Q�eh���\���?��Vy��:¨
l[���yܘ�.xR�P��L��ޥ�w�73w��Jk@ �lo��f�N	C�K��%���� {��S�������2:�~,8�N5�`��4!˼<��F�ÂUY1�D���B<k0!��������d"�"W8wS�$u#���Ύh��-^*����y�m�:G�� ����h��R>�V���׎�`U=�z���n�x�?�$8�\#��ly��h�m�������A2�2l��q��B����?�sb��K���D8�Z��3�T�;�V�.�X����q�{�~�aq������+�G�vv�Ұ�����F$����V4�X��L�b�x�*Na��H��s��l�L!�5�Y�CDCҗ%ی���͈�mqv��K�,#�3���F_(�F)��S�T	"��k�*+tu�r��f����(To�H%��j/�r��Qs.#�p;�ѥ�/�JO�cC	g+7,�'iС�#��2��]ܵP넶���>�x
���Tu���4�����>eV�	�!��@������[��~���J�o�S�A�_}�}��F�D��ǭw�5)x�ɡuP�(JU6����Fē���zy
m[�����������'n�ޏ�Q���1�W�|����R�dʳ's��Р�j�g�cF���|����gas4���6ėU!i����Fi��L&�v���C_�Vzm�o��]GS{%y�\tP\��L���
΍h���2�Z����hW���%��֞�zV�Qw��������%�Y6D���<�$%�M}�K��5�B������
�k��`�f��H���������#�M6�W*~!�LE0YP����/�qĬ)�e���0S�ÍR��>�˫��;ߊ�N�#���%'T1���y�^R5�Yz���,�.�|IM�6��DFCRx�M�BS�`&#��c�<�I+�~�Y������fo�J��(����uݪ�QK0㵝���Օ�����d`2pN|b�ӹS����$���W��å@ɾ�D��hA-��ְ��Z�X�˥���VyqB6�x���2�y��W3!�����Ν�c@�o�}��͐� \��y57��ز*�C���.uX+�MT.9�򣤝�^{�ӷw,M�����p��9c'�_�=q�*2��z�m&��V���X�? ��j�2��(�X�I˿I:^�hM���>��|$���A��Q�Pu�#<���
/T ��|��葝Z�z ����$���Xτ��9} %ݏ������
�{�*���O!����a����%U�ٜ���S�w�N�m��Ӥ���,�}m��lD!�T۳�e>�P�0iE��-�pQG*`���%ŏ�(��ej;�Mnhx�����K��Y�`C�� ��68����"�2�.B�!"`����z?�u�N�b�c2���	T���V���=�|���1[(�kA綠��t\�V��#�̑Y�*^ad��'^��`oOP
�����v��Iq��M�F�f�<�4�
N�&0j���C �:rCHNǀr�`�%k8^��7�Bs�A�@��)Ͷ�x�7GO?_������(yA�����8)�����P���cD���`nvJ�W]~�+10c%��7�n.�|�MA��;	�)����g��r�S��%���,�|��$� ��&_���3qm�ە67T�%KA���l�l"��mO%@ $Ow��ɺtas�yRPn�.*Q��?�����,�H6��ɤ�$5_tF.j5��X^n]�o�O�FP�OV���o%��(���>Q=O����fn���̮܌�Ѩ@�'�����po��k$M�atsǠ���8���]]�u���I�"��"�V#�E�˯��vh��q$#����mƹ�u%ċ�8<����<[�S|�@�z}H
��3p���AC�{׭=c��\�T������KR�/�[�i��Uu?�>�YD�u�r���K������-p���)��_Q���sr�N����]2[�;���b*
5��Ȉ�gx�s˿�	�5cz3����AGΡ����
������B�z�K��Q���5�Γ-VE]��v��u�m>��4��w�O?s�����n�}Rp�xQa��$����J�i���?����Yb+H�[�(88O�����3X#��?�d���� aAd��q���Ej(���,�C܏����?��@A�`�3�u.ב�v- �:}/d�.b<��d��@2*U����5;Dpa�1����t��lgǦ-�)1v5'��1@��i�fȤ�ZB��o!5,ޑ���/W������ZΎ_n��n�����0�v���-�,kmR���=��g�y?N¶}wZ���J�<�#gx�㼬�%�qh;�Z��e�6,�}E���ddb{�z��Y�v��N�*��I�����`��SH�Mǜ:-���EmM TZ��*������va�M��>�����j��@Iy������Zi�[�"e>B��bd;q�X6�Zr��[��[��F�\��p�"lʸ�>1*����ڈ������{Κ�@e�?��4(~�������mX!!�;�c�K���2��O֘��՗�=Z����8R��U��T�I�N�}���8�����3����^���^p���ƒ��/�c>��V��OEϕ� ��(��jwl�"e��)�C�:P>ͮy&ld2��O���;�}{�\O]/��6�D"MkL��1B��jVt�M��T�<M����#��MK�)�f�w����X��_ӫ.Xu4fj4�g�Qy���d�/��#
�٫�$bS��a-��[���D?9��l�_��`�g A�����2J��/�芣+��.M!���*R|���B�<�I�ĻVv�O/��Y���?�}3��!�$Ќ��9�H
�P����kA�|��!����V�P߶cXg�cE��a5j<�v`��VM�X/�ρAbJ9M�:�WX�Ab6u�2���Ӻ��k�'ߝҔ}��=���(��[C���>wV��(�	㴍�`I���K��lE���X5	&���-I�(��q�訽a�M��������V,$��{�y"�ic�hVn\qP���W)�ԁB��ɓT.�B��E	z��E_�)����S��r�����ǲ��f=�Vuq�L�Z|�`*H�S���Ukv�"��2I7�B9�n�yl2.���/�t��:���x��ױ ��r�4�L��'=�u���B��*�KI��@'u���g��]|����u��u0z(��yλЊ@�����IH��בT�6�h�3�����	'�a#�Kш��+�[�t����d��ΔD�u��p��:AQ��
PZ�M��ܔ̝�g����'Ẁ�#��=�>�C���)���/�4��~qN�PzR۰t�ӑ��*Lt�Bw�j�Q��[K��%Oms��p��0Rd�\�!_n�̀|�4�SG'^�5�,�oK˧�65v�1�{ U���f�;�#��z�r"`k���~���dh)l )��*��q+lkCD� l�� �A �E8��;xv�R��,��nb�fv��X^l�s|�b�0`%40�<�8�xy�t�����iӦ{÷~��7ޭK{�h�&��LB}��B
\�r��	u�'�a��,ա
$�5����\y�w]) bO�#�B@u9Z: >���'h�o��N��L�9\��~���{ќ����B>���T�#Q�;��+܃KsM��`֟���v����/&�䵧ԧ�s]��!rV�Q-+�.�Х�@�v`�"Ql.V2�������:���5,=����R������ȿDN�Y���7<i���
��T4�
���U�Z�"��X�#&�?�]@�}]|̐3t;�S��Y�h��u���y��-�@YZ+� .Y'c���F�$Յ�,$�5X�/m>o��y�D��]� ��$�*��|X���(t\�M��99���Y��O庮$؉�i���'-x����ЉN�k�Pt�F�$ L�j����q||�����r*^6W�\�!%0�@�i���ZKeE
�5ʆ�;�]���\��l	Q��������h0���K�T�H�g�[���T��;59	HAr|�� Dݽ0��V<�	��=ҳ�RA�W"�Pzi�w���|��k��v�GW���*H����W��������N�7���@�N��I)]�e���6�K�W*m�g4���S���U��-%X�F>����������d�PO�7A������T�:[�#���v6�+�QJC������FX�x%�]?1/xS*�8�\uz�/.k`�&��L8�k�pc�P���:��i#�,�WǬW�����L!jb$� �'�Z�����O���Bj�iW��[25kM�S��=G�����̞�:�H����g�b�J����Wua_���̙�}�� ���  ���o�%`](���  .�l2�d9�(���)��n�43�G~�*e`$�(]��X^���"*Z�#r��I�]
B,��+�B���b�H��O��T31pS�O��%�M7�#�)>�e�0�� �����F���c�.�Oj�
�֔}��.�-��5)~��I��?fj<�c��,�D:W�-�=.�l�x/ބ�� hu������hL�ڤ��JCξR|����J�>u��8�h1[�!�pr�>�i��>�`�2�}����D�%��6�R�H ��=�J�|D)��Wz���0�Zm4ձ���/FCa@�<���^�����n����� ��!�B��������R5�u<[*"?��S�ir'�ȝ��lkX�%g�zB�1)�ۻc��Z��d�L�[��W{w:�>��5��}e��t9^K�m�3W�������_���?�^e�EҘ�[enl0�{�l9 ���2%k�<S^���jm|�s��N9�-Lu;BZ;l���M�$� �АP���62�-@�’�{�.���"�=�&))�<Ue>��BB��3V���pE6�Y���pM�e�:V��Ag:9h��C-�r���Tk)y���\/"��B>����^4	i��Q�l�Y��dzrI�ŰU�	��[ݵ������'m;�C*�V��95ħ2�~��}	���0LG`ޤ��(��Pa��k&�y�IT>����P37 �ѝ�d��xuH��� ��<B��*jh=�d�_mZL�i�Ä�0��60�
�,D�lVd���y&8]��ZT=�Br55h�j�A�kN�"����5�`B������a6�1k��������\��J��ᓀ���"�##�]����7u��Κ���)�r���2YqY��m0	��A�a�^'��]u���1�g�i����Y �
���J�fr���o!����z���˦Re�ҡ��;�$�DRo)��	���0��M(�E����Ҳ3�@��c��~�
�g����Y
%�0�w��8Ώs���s�1���Q�̴}��!-AVCk����T�+�X���6�9 �D#�(e�a�G|g������b�DF����U��y)>���L�����|�RO�~�����0�s�%lv��I�����
7����j��$W04,��/+�0��6M^�5�o����|U�����4��m��^��*]�9�K�M��ؗ�=q�;���`�)��=�����{+�á�����F���wL?é�������!�����r���J�Bk��'+r�����&X9��;V�� �S��m?��EW�>��Y��m�>@T���>�����Lj����r�1LZ.�/�Ls3N���7J�-���`�(����x��K���4��D��3�'A�C��ՙ�'���R����K發V٥k���c�ҫo�v�jT\8�J��yY�3�$����~�q���2K���6E�ä�|
��:��Yl�� ���M�?!"��6]��{ɡ� u�"{�v�l�Kyd�IO�@���E�'�ۘ�{�����a�8��;MP�������bb`P����|�ƈ��Jm��
 ax�W�lR|��'7�Z$��G	�ra��L�}��h�x"\m����>��Ӵ��\:ws�B�@D��@�0�bM[F8���������ڋ�cXH`�c��ȚS\��<��`��@��v�9jg.T�����˖�ľ/?>���f�C��
إ|Я���G��,)e�EBQQ��[B3O�D3�y��ެ�@�k�z�n��G�&�Ū'�u��p͡���!7_W^�}W�J)Y�\b��W����
 ׎P��pw�P���"��ga�v%{0�d��th��k�)�2i<��BULM���S�*�i5�`_��X�nᓵ�������!C�@�����p����N�M8��˩��y�P�����sg6�I��ͧl8�w&2������3�n� W5�S7 z}�R�m�����x"�
��`�8ra����_�SX��W����9�'`Q�5���,G�����!-���I���i��M����/�i��2�29�����g��� w���j���w]vDl@S��~#I�\��Դ�#g��{e�e �zw\�q��ھrr6���8@.C���m��q3�0��05	�2�W�䇗�Q�^�`�$�W��l��u5[dA���.z�?�
�L.�4�V��%v�XpԂa,Su��{�I��Y�O|x��\%���(�͎-}�����s,f<Ǎi��x�PS�6�}�/��+J����]����y�����E� )k�����*%�_I/��e�>a�8���C#B/�㻭�. �x$1���\�v�Td�����������%r�z�����/��b��ob�Ư��@������>�k��W
�)�>�=MѾ;Z��C�`5S�~��X�ӷ5:̋�Fz�E���}���n�+*+@;{|I�@���d�}MP����p<�ʡ6C"�8� �Kx��h��[�N��é��e���蔚�����D�Uh��/�%�d�Y!3����ͫ�a��;���fR.
�
oK�+���8�e�FXg�:p�<n�mR�����U�dpQ� �t�"n70��]	�U�����Ж�S�'����w���zl�訔�>^�L��f+���^��L���oҎ����+���X,p#�kk��S5�%�d-)#.@�'{,��:c��	OI��:zYؘ�P��E�0����"m��?�.
�^ܼ)�vo�e$sE�hI���zK"�k�K̸Nغ�֖����4�L��&�u�O:M�@��sU3#"gJ'8�vG����0Q�~Q^uy�_��67q
�*ӈd=[���P-�>>Q�����w@��!�z��m�r-_���v�X�&�9�����['�nU_o]�.I��P{r�a�`tXi$�����P�8�L9� �����Fx�_�Ӏ�)(�����Ȣ�lہ��ͫa̚�~Hw�p '���oǆ���^y[�����A^��Y�2JMo���[���)iXVP�}��K!���x�W$� ՞WI&�)�7%�����dU&�X3&�FrW�co�-����jb��;q����Y�gnGZ|J[���g�����'2�X�(Жl��iPp�?K�/Y�^'t�:�9�뮞ض��(�c�e����\��uSM���%|�)����<(��ʭ#9¶�A˸�4��T��XRD����J�"�������5j��J������4N��d2s,)�3�b0�l�&�^�C/+E��<N"_�z�S����\�e�'!vBJX��ܫ���u��\���|�P��;�$�֒���jzb�Ȩ�U)qB�9�N�碜ۨ�_r�CS��7ީ�{[5���8O�����%-�WY��_u�Y[���N��(+�Yм;�c���;摩�^K�|g�92��#_S}��_�ڈ��(���G�����p�� ۃ�FV|?�r���3�wk�_�8�ާi�]��J��W�vup<�_}_e�SƹI�nE�x�D���k�8����w����*Ѱ~?p�I#n���)���΃�)�U�tPL����ٻy;%W����R��i�����f�K����D�?E����	���j���B ����� ��e�(ú�4OQ�b���G*��X�W�V��:���{z�BB�Oˀ�jMg�7ij��@��g�#�AFB�� �;n��V�^S���������i�aϷ�|�K��n���͇�H���<�8w�"��c�7aW�@����'{���.��2+�dT.�+�_4�&_�dkne/_� ���c��tʪ��(�c�䗣Qc��$c�9�SK��R�s%�8�RY3�R�yXXf�g8��R:^��D���<vW~�Ϧ;��8`��ND劸84*��t�c4�UzB4����	E��D�����$�d:U�p�s��kZ�X�u���Mtb*�)�6i����:���:U~�l@���d�<���� �4��\��\���x/�P ���*h��95o�x�Q�;���<֊|�d����G�Ksi���SXB{>	����p���M�
�K#e7,#�{�j��9_&��4H�\�s������?�%�4g鱬0�`�� x�L��ah4%���n{��,8�'�>�����^zCڝ�מ�&0�xa��Y�klSuP�τ^�l�b�n�K��UP��$���2�d�e�̽��&���*�+�C�e�A=�m��x�3�r��GI����؝e��ج��,>My��h�]�0�J~j�)0[h��͎���ge�X2������i��������ڧn p�x{Cӳp�]d�+�� L�(=��,�}�p�Zw�E� �~	0��n촩�b�Y�~l.CR�}��q;����d܅x SLumUP_���C��sY�r�hze�����7��\��-�k��&\�0;P�Ⱦ�ɲI�N�;�֞[@����ϡ�a����ص����v�L/�B7{;�D����!(��� ���ԉ�ML�j��]+�}��;��$f���T	dr�z8�@#�о煪����[�'a���A�Q����2���|�$^��ª����E��|����ւ�*��TQb�pH1*��r^eH��	�N�/�ӫj	�E�<��/�!Q����;�8�r�i΋�SE=�2����Tv{�iDBE��v#{q�2	
ؠ����t	1U���w�F�^��Y2	��F���v����!�6�� *TϽ�Rm6�Ҫ�C���O"+��K��rV�[�Oq���5
�
G#��� g��8$��`���.w�Tiv=0+f-kռ��=��Ǘ�"-��f?�=��v������Yz���b�.����b����݂8��!��'l/t�o����I\���}:�[uuI�z�� � 0��e��AF��|���y�]�f���v����e
0���`Q��K(z�������VDu�f�_Z�lR0��$���a�y�`�x��?�/`z�&-_x���#�K`��r"^�~� �ޮy�{�/���p�9/�"�v�.�a	���=~�����5s��ו}"nfӣ��~:�JKquW�jZ�铹t�}��"�U�Y�y��{R��`w<�����\�u����v�Ɩ�¦�CG֞d�����[�$�ypePc%������'�"��탷�s�LT��BrM�8�#��ߍ�En�GwY��k�k
�&_純�l-�AB�y�1�ڜWg_E��#x�
-U/���m1z��c�C��i�"GR��g`�/�ʩd���~W��P�S���6O%rR��C��"&]v�����S� +���a=]���6��9�eeT��>�=x(5 �#�	����c�~�h*T��1Z��epV��3ce�[t�Z����:Y1�8U�fb�^�ު�J^��_�&�mϿ��}�!4�V�2�DՈ173�5������*�'��J��N�"�2h4U>�]MRޮ���o����D�5��.8���.?p�����"��/9ٍ�ums�,�� �W0v�rU�^uxoZ�n�A�ڪ��}����P�a��䠁��Ր��$$0�햲�,
����ZC}����b�֤d�Er�a$gfG��}P7��V�#cjA��_��0S�L~���-����⛐9e�$���
���32A%�u4�Y��?��O���8�嵩��kH�Z����nt�1]���@���� �\��n5�V�'���;�5���.ȫ<T�c]��?���{Eڵ�ү�R�ٽ��� !��i���_��Da5��r�!�ly�Η���̀{�NX�<���]͘-��<���B�'�2�{]�J�����#�$��69�f��k�x����6�����$����7 {ڋ豤Fj��P{�FS��؛0���]{�m����|3˔8M ���LY�8,���B�9���[H����&����
L��\wV,�����7T�y��,�Q5J[�$+� ����HwqJ|	���(��<���6J^<yq�]%�l�7#�kv��}OkbHf�uze�(�O���!9���흦/���tÁ��OvC8�R+�͡z��h}�h��j�=��34�%{�!�lw��8�B��֖ ������+2=�T_{f� A�[� �@�& �B�*�i$9u�F�t�"�z�td���k�&�.��g���Wn��-�[
K^P.�IU���b�Z��>��lpz{���D���$��tU��ѐ�囯M�P����3�Ȇ��	�A��l�N�*���ۉ��g��B{O-���3�!�6mZԿs�|�"��͠�r?�d���B-��d�u��K�4M�_�����lpr�� �M�`���)J��Gk.��ٖ��5�ǘ�1{���OE��~�����V����Ey)E��{P6�7$��勶k��BgQ��h%������tr�$�
���iCA:U�]���E�O���u��Jk=�`ҼC��ަ�W(#�p[��w�+�`���Zʨ�>�����|�s`��&���Q!���|�`|�Ƴ.h�Ŷ�k�u�Hkj;�@F�w�Y�c�� �S�Ғ��#%����&�}o�;�D��>�<�})Yep���zR�� ?�@�����l.`���@�'��	��v��mҷ���F��v�S���b�ީ3a4F;7�^h�f"z���l��<��LK[�F�����/ ۈ���'�"
Ϳ��[{�?���@�:��;��~T9��A��Y��-�+���~��I�%��p��f��!�l㰅+"m����T��Br��bC8� !�(��7��@�b1��&Yݽ�,�H}B��I��C1@Gi����"ՓֲpR�����1!�rCC�	Ǉ�ku{�`ޓ*�N��J�i{'̹�c8��3�7S7G���*�m�K���Ƅ�BA���ˀ=��<t�N[�KT����u�*�ߠ��pSo+�,O�!�;�;dQ�ʕF,��i����<8
Q�!�8Zs�^�DE=��gT��S$��O�L��	R�<��rK�6��.а��(�����_�4�52e��1l6!�1��|��� ��  �]����D`{�ws���}
�ͪ��u^"�����͕)BhAB�e�Da)�N�>����@z��8A�I��b��8o�^��`�}NM2��z	�%��I(�*��[`�+E�aV�/�c�\-�#��t�����K��� A8��딪����!Tv]ȧa�#j�%,4`�6��W�R�c�L�<�,N�7hՄa�R���x|a���P����`�}� �C}�N�F�f���qS=���]�i��9���z���n���&Hy�/m嬥�Z�_"�� �ɺ7�6�Y�
K�3VԳ_�\"A8�� ��V�����������l��YK�f���2�p7��ڴ;�˅�����~��߱7�T-̲��J�	(=~�A,#樀3T��3�?��_�Ҩ��!�t���ܴ}P��d�o�L�0U���C�:ǥN��*}'�;����د��A?�:���Y��@�X���p� �$[��颉}j�-���ܯ��P�`����S2p�/53��'l����S����B[�w;�[�h$��)�n��=]"ܳ�A5k	���W$=����t՘r��PUG���AQ�U��:-���\~�� �za� �T�Ga�m�	k���K�C�J��V��S_?p�'�s2]��4=�sb� ���:_��a��c������*��6�XI�R~�(���G?��[��H\T�7R��X3H��� rE�|�c �׀��u� =E���Y�,>0	���a��ŧ��o�0λ��SD�qX�(;��7;f���6���IW�L4�u��A�-���?�`ӫ��lЭȚH�o���Pp���[7׳�.�0"��(�n7k�j����jB|s9ςF�#��F3ՄM���"�!L�V`��cI/~Ip��� a�����u:����J�j���u��Y�2�+����<P"�Eqo��N̯�u��%2�Q���f'wr�O����6�0,�oτ&*��@?�B���F�����4��i�'�0cd
 ���5�?`V�u����VO�g�S�h��ڿ����
\Wx���rE'AsЮ�tC	��
X;���]��Jd�G,���F�����)���6(�ǃ���D���O�}�c=�ǒ[g��w,��7H^���eVz����3��s����?M׉��n�'�:m�5��pΐ=�у������z��0��M�t&��W&�|�����^n�:U	��d���q�B��I���X��T���
��R`A�2�OIP��_9�v����V�G�	���eJ��9I��Ϙh�4�͡f����l�n�1�7�o$�H�U���ez�h-�+`�Wl� Sy$p"w,]���ϵA�V_;mռ�}+���疢�i��8;F:�� ����ew�[���Z覙�w�T��w��X��]��Ф��UZ\�����ϳ|��<�%�9x���3�J�n�����8B�toq+�a�G��/g���v�d����x�(��t4!�&n��b��n��m���B}�����\W�u|�;/
c�]eZ9\���3sK�JU2ĕC�-��dҕ�(���SGǖ�!��G��E-C�f�Ɋ�
(z.6������Q!����Ds<��S��v�q�n,�4(��g���4�#r���T�TJ�V�s�h:o���h��b�G!'��N��m(�_6*x���g�E0}�R���p,�z�$J��Cm�\m&����� o ݧBM'������#i֚50�	�,n<qB��?����#}���E){���,��Wht��%��3�"�|���c��������Dd�Z�������T0X'\-=��£���[
��]`���X	eKX2~Q��D��ܔ��9��"=� b�׎��}�)��Gªu�訳�R=U\��F���dK�pI(�IY������X�w~�7ѳ{M�'�ʥs~ڏy���Fv���J>��l5����	�Ri%Ά�-��"!o��\h禕p���qs�He���i����$8h����������ô���f�h%6E�"V3�!�E.�ӗT�s�%dS�`��Du31�G�:Um���W�~�j8�w�F��1]1�$���M/N����a�0�\D]��i��"�� "z�>�(�"��k2�������o��nlФ�t7�8�I��~�Ex|���"I�&<���?�́���h'g�i˳#�2�Zf�h��Z�K�z�~ϴ4�����D6X�OX:=<�F]&U�[��:�x��[`~<���l�b$
E� ���,������^��2ͫ���ˆ�hǏug�<�Q�3�z;����7{7������G5�,�D�j_ɠ���쁫/%�'�~> �m�4����.�a_0�ve�?����Y��F3*տ�(q+sN�;s!�9�=�  3Ȋ4ۉ\�ӝEx���W�Mj@����ج�V��]%��.GD�?��T-#<O)��q�?����a��a]�S�>���т�>
�����{�@��D�����R���~�̀�A��#i?�7>z�vgl��-
�����d��,�W^�����.o���JҔ@T«��§��.e�ֹ�{A<���5�0b,�[U�q������-�Q�H��> ��u�a�z�_�Br��%��\
��2��'�����Ϫ��e��}��~y�8��`���O4��j�(�p�2m��CΎ,�3��t���o����/2�Yk�b�i��#ĸ"��*��K?�����Rfi�l��m�]��h�������ɥ�W	-u��O���+��J�@;o�>��&�Q�
� ��=c3�AВ2|G�@a���^���x�(�P��i7�����}����l�ֱ.~�|�6�ۉ��|֯S
Id��.Rp��f��r=�7>��K��a��x���?Ƕ��٨�E|�⾳� (�=�;�;GgG?� Q䷂�2"������{T u�фF�I��>�����󕡧��E4��q���\R�K���B��6�6Kǯi���'K?��PFg�*Kb+B#*��;�����՛��S�����_�T�č�l��B��w��Nx�����Qg�3g��|�:mo��)�6�l�͌�����<�߆)W��S��]�Y��� �^�p�sp:7�0��m|���ĳ�>�V�8�3c<їA�8z��?
C)"-?�_
�i�iL��}��5���RJ��є�jKP�5��oL��3,���|1�f�.��v	�*֜�3J���kTpr�)0�F�Dr������sg�%s"�%f6��o���h�ڷ���[R�Ŭ�Ɋ3��
��g��g����r�+�^r��C�N�-SQȟ,~����d(�R��
���~n�~C��kn�ր1~�������nyw�*��{'�3@�*W�D��=���2c����m�D���=DUQɗ���C��Hwk]��� \eQ��G�����Mg5]��l@� �8oB ��&Xg�`��;������S�����᫏HT����l��X|Þ�q��0<ؘP���}EO�1E븫X�pY;̺�>�wvNn����Kqk����hQH�1$m'%���]{?u�қ�B�R�e�H��ۢ���D�A�LG���R4��Y,q����k�}�k<�f$"��B2Y�	cP��d�Q,B�.�b���T-w�q
O��'Tx���:��f'_�xMp�l��F����>?�g�7"�y�.��~���(<u�ߵ�c��"D�#<�a�m	y�1G�� `�k�]��|�q�'4��1'P�. �j�K����݊�8����ƇdN��
a�_:C�`��ߑ�
q��.�'}��?}s/��˝˱�|�E�����s����V�覊-k�d4�8�Bnײ4��3����;��ƾ���וWT���¤9b ��{�#l}Wf����{�DH��Q�M5M�ɄqT;՝����{�}�*�о���rR����&/̐���v"��f�q��uN�H�p��.Fڙy�1��Nj��O��8�?���M�����P1	�@��}�!�N�J���#�9��E��@�6T��B���8��f
ZrN�ֺ|��	�Y��z�J����ߦ��K��]��t&������Z�M�ul�p�K�~��--rꁴ��B�z����O�U+�yůx�$���m�kYj}�@N��  �]����$T�����WՈ7)�r���+�|��FdJg����ԁ7M� �9�Y$|L���#���f�k��D~&�ت��z�D"fl�F,|V#�@����7SUjP��_�7I��oi-<%Zu�#���N{��P�M�OJ9��P"��>���cBj�z�E�BȔ�U�w-��e�P�:D��\�X5@�P ���ͬ�rm����a8��C��D����n���/���|��2礉����2�AJ{@��F��Y�CM����۷	T�4@i�ҕ!�t���3-��BlJ� z�,_�Z��}�_|�����5�u�	/`������?�t��J�AO��̧�&k5�>����sg`����g�A��%�����hJ��x8�e}�S�ۖIƬ���q�$7ǌ�5ݶ�JeC)n��aP���Y%y3`���1{U��U�0�&��coa�N:yr	���	���4.jQ�0�՚�h�����kz/6�����מ۩��i��5��#5 	~��Pn��F�L@<q�%����#���(`�6h�A-�%�E!��<l���C�+�j�_N���կ��E���f��ƅ�q��C�������<��Нq��	M��ӽ|w��,5�A��\���\����`r�?�������Ɖ����H��i�xs�J��8�fnz\b�e�u��xчO[�G��u�Ƃ���7��Jo\� gJ���
O]�\��8e�[��+�d�T�PT@�:�$��xё������8�>��V�d��A�w,�+��g���5��5࿡
��uxi�a�?!BAcj0vy����E7�����/� �`�����).�J��1���W�u(����|]�~n�f�\߫]UҶ}��=�?�M������z4�M��h��
�����������I��ŝ�05��/�:8Z�<f�E>���*�W��23<	�YTT�8%0��(��(��p�z�f��(��9ve���E����[KJz����zSd �wL�*���O�|�^lr^�j(c��ø^��Gvߡ٥7Ґ��7��&�rx� �əv��:��r�Ҫu2�l��*��754�N�L���$h��]+�gٵ��#�O�)J����sW�gM[� l��d�D�8�o]a�'��i<������D�Ȧ�υݝn���闞����:Da�$�G$go��"s��h��<�Yb2\WDZt�l�:��m�~7���a̃k���@�Ռ��X����h���a-tk�r9�l
��7��Kp�;q�CYx�ۦ�������!�8�{O$��<��ΦO�5�J�%<�ܽx�!�/�W
�gl%-ؠ�'���aG��q��8+T�$��%�8]�r�N���Ƕ��>+��:T�Ŏ��ܠ�P.����V8���7�f�W��ҝ�Ĺ�W�����=��ƚ��Cr�'l��!�q�E�m��oM��U����`�6����KaV�E�?	�����Sݴ6Z0&o�'�)��؇������2���HC6(>+[�
�K�~�22���~2]Z�!�u���y��0�4j�)��zv��-��͎��z����|��e���zD�<�t>��5�� Wt֪s�Ʒ?m�m��joqdMnR��e�tD#u�x�=���2���O���w��n��p��o��jNG�]t��}\3���{�w�����WQO��|���!b,��i�Pj����ا���7�H��F�)�[F��>�g�֎�Ic��bj���v[)^6��4�9�2b̔[v+���sRR���l���c�A|afz������%f=��R�qx`�� $��;��W�������N����{)cu4��:��I0V߼�X�s!��s��^��=����3��TX��	��Jy}p˔|2�/f(�l�0��/�W)=���^��r�(Ĝm1�`�$%��4�k�VA �K����i.�GJMSé�b�0x�U��Jv�ᚍ�����;�:��QW�Q](Q�YlC֪n���� ���}g4F*eD�p��"ӊf��V\XS��k�Z~�����j��^o|2�� XׂY8�m�����	+C�䫵�*�Ok)2.�'��k hik�6ї\��j��+嫿�bX�3�3������`�s�����gZV>4d]pୌ��.6�����4?P��=�W���v�@�8Un�Y���<����UL��MxZ<�
˜��복�þ���v ��^��ء��^����S�kࠆ� �g	g�j���H�q~��$�zaa?�Xb=���ȺlI �&B;�mA��]���\���;"t�;��>�xS"�#s5F{�nB=!ބh&6yL�r:O?����l�/U��.�Q�|��8��
� ��*f�>&��&W4֊&�6�M�ë�W�.h����Ī˄,s��ڢ��O�v�d[�O3��g��œ�;�Y�<=������W�	9�4���P�&��-��i�5��[��FQ%W��0�E�����%G��<^l��,�}��~z��UM�	�Vw�O�X�Z�����Y�61TٽiL��D�L���˩|M�.N��"nC��AƑ_e_~ �KQ(��̨��{��Z%�k���k����pX��浉��)E}0A��y����;�Pq����i�{PQZ��?�ucxG�\�N]%�ysjM������LO���ڎ�Xp�:&s!��Y�9ȉ$t,(����n��M�d����8G���ʴ�,m�k��}��A*_>{���J:3�E3˷%���f��'t�Z*w�<���������T �S�j8��ς�G�I��	7$�<��ˠ�ZjQu��+7��P6�?�Q��Á^�W���{�ll�*{��q�j��S���#v�Q��#��<g�X_U'�J���Y]�Gݵ܉�]��1nNx�؂�Az�����	]�6�n���F-2�LF"��j�������A���K�]2�S��[ ���$�!�b�U1'����삲D����������^�OF�ggy-�;�e���Q٬4B4�"��e��sv2���;��T��L�-�ʩ$/�K���f�C�4�����z;�����åH��jq5���BLהd.kj �h4�|��f��D"���{�!B�h�"�O�^7+�r�u�+�џ�o+ܚ��YeL�y�z��LM�a<!e&}=e��ȴfo�v<ـP��c�/���Ġ%������	�~��u��Yi;fa/Ms`��,L��*����rr����o�9��T`Olm�j�����%���Us����D�6��ַ;ӆ�:��Β�vh'���e|�nՖ���qi''3�َ��T����[oĿ$�h:�����̱�FT�*vb��,����|�]t�T���8\�'��ӯ�b�_��8�)�b�����І�;}���B4���Č�L�Ĳ0��=��鮣дx�Z�i	AE%T����]3!��I�6:�>q��s�"t���<0��+�����M�� �#�k�iye"r��?�|,�)�+q���>6���U�܃l�����N�٘��\]�����Vl��4'����eԎ�훱w��tR{�y(��J�.� �Q�T"�;EI��c�Ps:��(���K�)�h�0�z�����=籍H�!ޅEM9z�#�ED�X��>�����뇍WGT��=*җe�fɶ�g���㜮��^�Y-��";1T��Cp\B�*Ƽ �b!���i�@�����U
�$]|�W�l��"֯O���nJ��Ua�N�u��3��e&��tk�䪅���.�<��M�F��ց�H|d't=�c*����ua���&Ա��P�Ǻ%��v}�� ��s��~p
8�i��ը 
I\�:lw%Tmc��̬ȼ+�.���b�+X@6�������Wf{U ���2���g"FI��8M�e�O�7�eTڿ�]�ZEv%�h��>'��j���\�Rh��݅�<#��bը�s��§������Б������e��~W�E�{6�/R�^'��V�����0dY��s�1��Ɠ41r>��ty�0��.ٱ��VY�U%UC|c��M͉^��:G!{N՛b��J�u�����Z22{m��q��4Yw>lf�V�c%������� �<��_��°��'HxK����w�.���k�	k���A����783��4��5�飵{�³G��A��4�o�B�:�����?��0����6,k&E�U�dk���lG��"�r��P�6�+|O�d�n;��<�Wd��;�^�<�C���s6אc0��Ǳ��0�����׳9���H���t`��O�ؕ�@�����2��X���'v�|�f�� W�&�����L�&��L�3p�۵Vާ�AS�q��1���'\+i]jm�~�t��g<�J>uA�p�T�V@Ψw�q ΍�q�p.���&P��nq΋ˊ8�tV�j�ڊ�bF^J���^�
/��5=�k��8�;�}n]�W�l����;��S�2'ĠY���t��r��(M^��1��/����l߭&�)�;-'�@XK����_��~�G���[7G�M�r%[ӵ^FF�J�v���" �#�1��*䘗j���c����]ge'o��L���\S�js�x{�P�s�,2W��V�f?����wK4��3%�N��S�_i.4�X�"�������m~��H6�5d��O�Ccm��f�1���A�8�o�y�3<�v���B=a�կ�u�@k"9��cjA�WU�hl-_ɧ(�_�K��|������9���⺲���:�μ2����X3�Eg��t��i�����B�e��`�^2���)�����	���֤H�!�Y�<Ü_�-D��vs?-h��0��V�Ǚ���e�E~���,�Gl��{�-7��׫��-��:²EԸˋ_��ڈ�Q�6n]����h)���b���Ѿ��p�܉�MXQe����Uװ(������0�e��c#n%0yN�c�%Z��\_wՂ�]����؇Œ�A�<(��z̤kPp����;����-NO���-�󰎜�Uӝ�CE^N\h���(ڑʹz���})�4W�p��|�]JP���G-�y����4U����GE�R3��(BT��T��غμ��ȣ�j7�W�.�d0Ŏ��D����N�T8M���j5���2z6�3c�Rd���=2@�,R�ϵGYSMm�=0�L�}�PC^��������Qd���rb�-�9+�qZ��&���q���{���eV��7 �QG3-�b��W�J��	��A�m������\������]�>=��L� ����4I1�L4��G�+�6�=Y���.sQ+�����g�A
N:��QWL��.�f� m�����E0��`)��o�!�}N���� G~��/:a�3w�/�g��v��6_��0�07fo�jr�	�|4q��`�Ť��P�.�Y
�4KT��=N����1����n6r���j���7ʲ-N["%��#��>���J���{O����OxN��!XƖ_ȗ���#�]��U�Oj�w��k�S�aE�f��vEʫC�l+�nD Ƭ�Ԕ0������/fA�鵓c?Z
���z��?�J����]VG�J��R5??��'�\��/?����g�<�xB�����2?^��Ȓ6&g;��G̴�#3ٽ��L�o�a����uEH,va�����v�����@�p��|��%hI�]G�ݸ�A>Q������¥��Hn���X#\�O:�t�e�����{}�f��9T�jf�K��~"���!V�-�W��͹�v���N/��?�ό=��p9�ڭ��5�WZ�H�D�y�Y��Ɗܡ��r�Z>mÓD���~m��{c>�.�����w��W!�-���n�@��ِ�_<�7���N��me�J����ݜ6�>g���Wfa���@�&�F�&�$�Y�5*9!��Tp�ly �)�vbx���x�j'������/����]*$�$�"=o��^.�����_��`�JL!P;��4�*w�G�i�q���D��-c����6��:�l�@)�@c��c7�#Y�9����Ɍ3�]�?E6=G����Ɖ�{Q`z��y渳�w�n��,1�������(���Ӊ�~�M��p����&5���s,N�O�+_[E�O"o�^��3��Դ]����"��L�5 ]G��Ea�ɗ��C�ջ�t��(��w;�G+�j8�f���ˢe�c�%�m(�G�f�����d56m&���zm��L����C���s��ܟ�=� ^1*+p�����	��U�)ݦ1{;��T	�N�:���(�>6�n�C?����C������Mb�+߰�)�8�%�x��{�m
p*�
�چ�W!�޻!Mk�s�Y���3��߽��:h˗���P:�=z�k/9��iA�6M(at5�p�=�f�EQ��Uۜ�E�az(��c�4���U��3)��	,�����h`ԝFoT��_�,n�MxJ� �y��,�pDI1bG��$�̼5!�VBWh�Ïa���2�˹$L��Z�l���a��t�%�HEO��9����./���ҖL�|�f���K�C%W�uLCW���2�&�8�QE	鱰^P_B��<M�wjy?z�����x�P#����2�)$���g��7g�\qRW�p��G;�R@-��%�w�:8]0�p{���F�����ѳʤ�,B�;w"���a��$�w�Gw��/�"���&����z�b�*�w�`��ۛWi��=&��E4S�f��3��%�U0�Z+9-c�i��O2���ȥh-ͤ�{�)�gq��8�Ȉ�B�
k�W��eK���.�&'EE�� K�WS�iFӆ�I��l70��F/����2��7͑�Oiڢ']f�}�prI��0������ ����ͷuB���/n`�@�$jS�],j*��mkU6	����_T*�(G�T<x�x��1��F�_5�$��;�cؒ����W�Ab̓�02��#��\:!�M ����[����P��?���$%��$������E���av��q��L���V�rMU'Oo�~�鎼&0��#�{@n��51��� �XT.߲50��DH,OÏYr�E!����A)ej�)-@�w��/��8��|9�`��!�#ؐp�A�ј���l����Wr`/c�f�og�j�
ﶫH[F�J7��,�x�Q��취x�(�>�ʌ{���n~c�=1��=Tw5�9���/xފ����ɲm���{z2����
c���w���6\�������`�-8�;����Th���`2_�3��6����!"d��kq�����R�^C��E�p��,)l������66��m� �G��Y��g��^���,}���z.��5�a`7�)���y�I�6V�i@��`Bs�V���U\I�l�a�\�ʝ�7�������*�0���b��X��=0�ڳdE����1P��.��@QЊ�Z07���Gg'Lk¤����~+����sA��G�
�p����മWs_���M|,���a���TA�A^.��R���X����:z��-ܷ�R��'���+�t��3�k�N)0�M�	����w�F�9�:hU4��C��絖\8ۺj�� ��R4���Ԯ�(���-�M!����T�߀�RFÒ�:t��NG�@�q$e�`�6�/z#��P#֢M������Z�1�SSfjl��"$��P��-��
�C����Q�pG��Q��타�Pu�����G��v��%]$-�����(`����yw|<+,ÀL�!��l�VsksW���Yty*�M�����#��|�D�ҰA�hd����������}��� Rt�r��F��
?��*�T��s-�;����ղf�&_h.�W�
�u�7�4�@��ք�֣��~?7���d��TΌniմŢatC���A|?gĆR�|";x)����Hڸ�"Z�����L�>_BT���c<ߑz=0��Lb�{H��l�!�1P�--�?��j��ND͋S�o� ���
�SX-J	�
�L��u��鳮88Vӄ�$C&�n�216�P|��-���f5Ҹ��t����.l����c��v�d5�e
5�&g(!4��Y~a��L6�L��d���@�ty�d57L��P<G�t��zI�T��8{2$�xoZ�Y�76o��_-�Qa"$�^jCR�A|HF`"�T�P��ss�7��#?ߟ��}�!��g#�h������C⇰���"{��y���s7��h��)��G�&��c�觧#y�0N��K��kU��i%���hf��H�l!R
d���uJ��|&4�S'V������(HǕ;�K��~S;a�Σ蜏�M���%.��>m��E��M;ћG�.t�V�6����e�[�H9=��̓OoصfӠ�c��&���m��G�>7$��.�BNix:�|r]�Q����v%��5�֝q_�c�f}�;}�g|��	�����a
��f� 4�9�圆��� B"�� �/w�Df�W4����m��`0+C�U�b񭥩��]����C�X����@���\����z���.E�[jj�	�8*�x(�KEt���oI�㶝����|R��]v������F�/��¸��I�d�]�n1U��{��lI~�����s3\,@��A��9���mءնo摶��4�hin��x�x4tWsm �2v�<�]tG�,Z��|��Q�	£�40���,��o�u�fk�~t�%g�8�����d��|�q�����W�����wڎ�:�����Ef	Z���ҳ��;]�CnK�5Jc��V_�#.�)Vfi�&'�P������,����s
:�F����,X�߱ԥP��N���"�v[�C��)��{��4�g�m
g�o�	��l<ω�|K6Nө�� �/�e���h�ο�5E�ӟ��`�m����6�6�K�B|T�s^7.��A\�4����\�<����zs+lD[)�Y8���F�Y�9���Jm�#Q�IwK�1:��nT�0N.���x0�)����h�]�j�kV�5�-��	��M��.(�ka2^{(� ���Y�'c��}�;�����X:� �N��Up~��u�&S����H�>���R���}�;v�LH�q�U���R��J�4.�[���k9�Qm�\�G�� ���r%HT�d�:��+�>P4��~��YA���8h�\��
AY�ĽH�/a(����������i]4d���[N}{ѳ�8X�<c>�΂9���
�Qz���]�H-(ks���Z<qB�� ��gTw��
��9F�f���9T���v����̶' ���§�XY�	P�]G��c�O��*1�����>��拆�w(��Xq��r�j��D��]	GFW�qx�M[dg�R�EbZam�5���1���VY���I�Y����r��T�O�tW�4��3����<���*��ֆ@�<~ϼ\ q���b����\j��yGo�����#���_Z�z\la��p��b)ǵ��5C�չ�:�ؙ㣯l�^s9'%U#l���C�#���E<������XU�b�z/š���R#��8�7�'�Z�-H�㤩�]	$r%�<������s����.Vtm�nBi6�>�6m�T#(�i��O�:{�LB�4A2ͥ��֟5�&���!y��I�����G�S/�eP�Rw�c�n��>�X�Ќ��j��7����T�w��LK��_]� p�h9��q��y�cX솢 ~������N��qi5M+���\^��$"�A�K!�so�^�q���������������q���h�o�H�>�Y��E���VNMjTzj�jH�ԑ!efVX~a"�X"B��!��
�oFC"Gho��J�ނ�[��@S�.�)\�<d����ܕ�dY	�U�F1-bF���|c%wx�y%�u�ek�&Vso��7�G�y,~7��{oL���mP����װ$o����]�ъiRD�d�Kh�B���鿣�s`�PE�#iI+��s������!xW�A�ҏ��g��1%(Ui
�=,�j�6��"zWX3߃����NO$NX`a�٢
S���R�{a�]"� ��u�=�72pB}r��� ���������N�.�����z�s���O�0(@�3F�r�'*�ƍ��c���>��ކ���K,�f%�D3�BZg�8j�<�NF�b�k�`�������ך�/?�����Hu�,�l��%�c i94�)#��/���|m/~$��M/=�>�ki��|�wkj�S
N����,�N(�*�KXtJQY��{�L���:��c�s�.��J�c6�~�i3O���5^�N�q�� �9�N>�d6�� wX-����*<�$��G�M����i�8W�.2�XG����6�9D6JTQ�@ ��4��:�L�+!qg?��O('�«�/1�_vT�v��__R����D�̖�fH`ٜ��)��2=��]U�����UB&�A�%a+�l^!�՛��W��R�eLzfx�2C��:pJ7�j���綸%Z��(b�0'���{�ן>+�$낟IB.��I�� �.�1�t�ߔ �1�N�Y��'�%�$X�i�/���:\�-���S��-.w��T��;ݥ�3���{6R�3q�BJ����@{��+~�s�o���7�@�N�.�Vk�f�w�U�c
�����E�qLY	s�M���[T�8��#Z�T^�O^�*��pz�&��]$�l����PQ+{�V؁�K�i=ԭ)��$|_��>@>���l���X@�(7�T*�9�`O�NU��U3S?�`G�%�dH��k2���=/�ؙ��X+�L��V�@���U�!k~��M�v9z��ʧ�W��� YNb����
�m)tDǯܨ�����^p�J2�[ܯ�%4�O����}˯�ǿMG�{�ƀ(5�����'gä8}����s��h?p6�s��c��;�ZS��%�&��ʝ:D�֐l3g��=�9�nK��Ѽ��vq��RJ;���o��sK���
�J�O��������;�N r%o�i�zH�(==�,���Y�7+�����i��ɯ6�D� (�:���@[p�5l�W�'�:_pNq�W��(�Z��F�O%8�x'9��(O���QV�Z�ܸ�,��g�p�N5����W^k�!�A㩩e^!Y)iv�UC����$.Ko~��-��J�V[>􊩲nu�x�٣�MK�*X��m#4M8�R��Ӏ��9�3�� �%�|P�ÎDD�:stv�WBgp4��U.}�+�M�#C@s�7l__#��n�=����0SQ�y�un��f�})V0�|Fi����z�%��7�AY� �Ag!�^�����#y��hb��g�i=�^ā�L�6QD�,Fn�Ǝ�1���da���v�!�骞-(���(���-;&7�uU�����HtUg��>�}�^+�_]ވlFṸ�wk S;C�q.1sn.�2Uh:�ΥEf�7�Nb�ιi�{�!���/�z�5����2q��z]�e������ļ{���:����ϫ$D�%���2�XH�K����
���Ly}:nN�ݘ]J�%��s�����$ɇ^.�0\��ߌ��&)�a�v��6�����Xү"�'���R���Xu��P��X7�o������-^��8��J�I�l8}	����j�JJ�*�+/��O�q1�IKп���&F�ˮh��x���{Z�=-?3� i'�
V���	�Ik�3r�ܣ~�Ԥ��8ݭ2~^�y�@����WydG[�
AD��)D���!�7U#zi9~c�u�z.��oR#֮d��3#f�G�h�)_{O��+�0I��*�Xyk�yoMQ��׏^���M����"��ϊ���(Q�����n�	���zvS7sԛ/��b]k���p����k}o:���E6��{Rf�䰝u�8!�e�Z�ru�����	��Y���!_}[;�s�����5�;�M L���Ͽ�h��X����!u�UT]/�nE'���U:z�k�1���\��bd@�+E�Sxȧ{u����E���*L��jQI\�zd鷃�ND��FQ�5�__�[�D�_:K�Ṃi��=ݐ��V.b�[
����m�k��|�- f�kz�Q==i�/O��Sm$B'��_�����2��d��[����T�+�E������x��;�
��䖚n���}��l�tJ KQ�Y\Q�4ol2*`��؅�_2h�a��-FS5�����n��U>f���˹��s��Q�h�5�������.�0Ek������ ������5��E _|�iߩ�SEs��f��`�\�#۟�#`u
%M��6����r�뙷�z���'�k`g	���F'4�1,�ΡZ"��O�}b#���៸�S�l��_�*�|�t�3���]�췯�û��5�+KC���+��RU��O�%��AUUt�E��;o~j�t�K�����z�/܂M��.�K�;sP�++�9.�
E�D �sdFk k�t��4ocx��Cۆ1�&"�z\lz(\h�Эn?��w����ncc�D�k��͞�w���㏁&��0���D�	J� Aؔćj#����Z1��LX,Ħ��XIA��CG{I�=:���ަ����]`�'kB;qds9��O�#.�=�JK(.F"�E�O���ޯ���_���?�ϫm0ġ�|_��K��Crp`ɉQ�*��Ks6+�
�M<�T"���GÕ���Qt�� ���j�g� �6�S:_��o�$v㭽���iw�b���Y��
��Ko���lTN$��M�Q��K�F2i{%Tb�	� ��J��ϖ+�ݟ�����r�x˧�)cM��.�@�]���w1�N����8���o�9�Rǐ�� ����l��h�~�t�_���ܱ78�;��]��1j@4{�ȞP�g쌵-u���v,k�8B��|d�V���[Ҝ�{=N#�� ä6~w#۵�d">ję�;o^��k����C&h{�%>��d��=�9�]
*8�մr�G���j�v�>��(|�
ޕ���
[4�]of{�O��p�����ŏ)�me!!*�R��XK$����ښ��\y��û�����ΣX�;?�.�����Aq�M�RՃ��fX/��=�|$Qn«�R���y �H*uq�ާT<��\P��vCx�z\�ɬ�Sl��IX��84	���3Xq�@��1XxZ��%6gi�nQ?Q����8���a���kZEde,��
0�Z��y�0q@$���[Gߙ��օ�M@�\ar"�B8x��������F�r��o���Iԁ���z���d˟��Ǜ:�ʎ���8�`�[�c���6M����Y��Y@cM�W�����")�Ȥ<t^��X��sW(/x+E/�f�{ͺ�_���	>�)��}o+Vd����sn�3J��@��D13+릈��ꠑ��g���/�f��"|C�L({N�{%z�<76`w����&�,~�S�����\*WJO�,"mHco�]^���|+�YPh���/�$�a^ɾ`ڜ�i6xW�?R&�F�.F�8�f7�
��A�=$'W�pK��`y���Ψ�'�K��{�"���6�[ �P��c54��)*�e}�NTԹ�{'i̤a���pa�7��+��F�ĭX�gp�qԹ��2��q�\�q�u�Zcr�i�x�D軋t^Ղ9� ���>��3oH<���Bw�l�"O���p� �vrw�*,Nˡ��C����p3՛�P���C��"_��U��:!;��4��cu0	�)�*nx�HM��<�1h�����ߩՈ��@s  z��J��E�FmL�f��Q@���Om&�,�C�5��ZP"4Ź�4����-8d��Rl5�o�ɔB6��Rs �H��mi����S��T��\Q�L��7��p�f'��x^`�s�T��m�(��Ip�L�7��u6�Q�`��3mk6���U"���Hw.y����	�A���Z����,`����4���	�wA��| �����̻!�>d�I�b���ų���#��ރSX�R
�� �
<׉k)�}���c�_��d��D�%6ڱ �p����צMgMZ�W)3:g}�[�䙖����D�W�q'4\CCX��bQ@|���U�u�kTl7gV�ںM��(�V����ww�5$o�J��+������1����?���XW�	щ �k��;�u���#2�ˑʑ���-6���b<�[��)J1���j�,���	�zΣ�eO�R��n�*�ˇ0!�;wM���J�uџP4���	��F<���n���Z��&O�Ɣ�22ʇ �9�:�j�!ӌ9?V[�D�A���
���"�N$�x`�x%ک�H;m)�r7��&[o�A�6���ۇ�ӣ��Hy(z�>V�����:a'�h-�)_ot0XKk=���b'�}]��[�B�l� �xXWZe�a%�28�sB?��j��22���T]QvԳ��y��ipYkt���C�����H��7��}o��P��u���ɠ�F�u���ׅC['gwdi�xA��"���ke:��2��Ө��[����*�KA-9��4�������;Ξ�5$\K";��~�k�ɕu���h�V�GF[8�y���p�X+o^N4{�t��@���j�	�D:u{,T7"���]�~S#b]�wSЦ[�<��}"��4Pl��T=]��J2�����u;9#���,��U(��j�mW��"��`C�]���Ycc��1�ɝߒ��Kbm�ǣ�٩�9�v�@���H�lUB��<��~��m5�%�Ѿ?���{���؜#���kK47�Po���ڳ���j�,��sDX��F��Ay6��`eau���ΰ�ß%��$����UC�7ÅEoZ����}��УK�9����ݜ��/K�K�Ǽ���~������Ў[��ȇX�����'�Mǰ xV]�\��0�| 1��)j�\6�����U�£c*��|��`�0g�9�mu�� ]�x�1�v��9�	�����Jg@~��4<�Bo#C�P������Ş�Q7��9Ѕ�	]xb�9v�:X�r���dkh}9��|}���=j<6���c��p{y��"Jb��j�V�3����M�2l���)�b�4|����NLy'Q4��P	��
���w��2v�G|����z�參+��ߋړ_L\��f8p�.Ki���DZ��2rW��>�8��:�M���W)�	�h>Cg���Zpen�V�2&�������g�d��q`��j=�R�B��5����Ő�ɖ$��*��8 ���^]��9���b����m�?���|������X�S��T�m'�p��L��w$rf�l������K���M��A'(e�r�Ųi��T�K�BXSVaG�p����k�/p�ϑ� ����h�H��Z�!�1X��-�����b
�To�)<*يv��3DXCR^|-��W�?��C�� ��TK'��|:W{��+�*U:����U�%Oh-��qo$��˔i� �pU�.�S���]>�	S�Ɣ��NH��}Y�L��;b"�73I]ؾ���!���T�O�rҶc9��ܣ*��c%��-�o��y��7lg"�
T�I�r&�g~D��/�GMN�oMu��n?����stW��oՌ%���Bn��&0��`��1{�zd�#�*ab����ӑ��t��O�@��k��P�h��X_찹"�^d9H_r	q>�aӑZVd�W ���d��L�������,�Z����ܢ�v4Î�z�'�N�r�_P����ҝ^*��ԗ|�Z�:M�<5�9s��L~�0}%�����Q[�1��t��B��Lm}P*�W�^mjxL���<��Y/>!f���d�P�ڹ���N�H�$ի�X��_��@H"�$+��Z��[g�`&:��B�iܭ⽩�Z�Q�}���ps_x+�i`�Ҭ2�(��~�L�`SW�P�?�Z�%�Г<�zw)�T��>�P4q���A--�!i���B������m�.����_z�@��(�;���pI��1D��0x̭Y\��t�G5%~H���V7�O��2^��~B �>�(�բO�Ԩl�6���<���g�6�)�d�I3U� T�(�'E8��CT��>Z�l+#��B1�Ï��S�d���#Ă�Y��uI
�I�R�F�M;�  ��c�[��{�+��*���!$��ǧb]y�5ȚɠkbO��W 3eXK��B�(z����("�4Q��M�V�G$�Vj>�/]"�|z�Yx?�{� �l�K�;���?&�"`(ӣR�6�G� �W�� �z�y,A�����/e��rL�n����8�'�Sf0��a�+	���62�-3{x*�� �'����+ÿLk�g��V�����R������uA8V��t[��8G��ӧ�E���\��b�>]V&o�{�S�'Ĩ�Pu�� ���8cg����y
�ȁt褬i�\��8$8�y	���p�Qn�ˎe���^v�D^�w]�iᆰ��;z�\�&�EL~�>E%g����u ͬ%����0c#D��4"���?��V�{eK�Хa(�j�+G��c/N' ۉ��҃Zt��E�K���:��t�3���'3Hw\O�Ytq/펢�t���F�"��`������E&���b\����أ��Rs����s�,�~z���r�x��{26X�֟�G�CA�T��=��h{)����;��5f+-U̴��L2%�* �4�P{�:C=�>�C���{V�h�|�_�V��k�@qVΙ�
*q�+΅�fz�cR��)%LQ���yw.Ӓ#&�rI�j�kܦ ����Gl��B�������O�$�]���s�t���H\8ײ��n��(��Ň�-λ����׉��P:&�Qpz��]WbB�G���Xu*���2��^�/�|�Ȧy����w������۳O����Hދ�~K�p�g�v����?�aK{Ov�PR �l2�ۅ���q�����8墳D��xlu1?vޑ-c�t�U����t��	�6#5�{���"�ˤ��\��i�e����Bfʕ.�J���G����W<�������y�*S�{�8�_�ۆ$�P�s��ĸ�ޑ�%�>j�6�8��T��ĳH���`�4��f>�����X�DQ�}t\�pGղG^�~���u�`���g�#fG+>��T<�'�O��D`���ە�yBM��:��N�+uE0��	o��%1>%���q]�(�o��m�uɋ绪���AKzˬ���I�ɍ�}a{��#�j6�z�c
�#����r�r���/B0U�$Z���Ƴ��=W�C�~�qak�[ˁ��Z����3)�}棾�� 7VP�xî��c熺����@�������� Ŭ�ܭ��� �_L��hc#lk���%���2���J����4�y��86N�m�%$�[<��d�hM�<���x#o�#�1S�Z��̫Hox�,�h���d��b����_ru��5�hlk���x4��`�G������Y}ORn�5;v��.r�s��lEsu���(�����k���۳�gܑ�����N�C/�6NS���nm�n��1
3�l�G-�6TSV.�'�`�ಁv=�P��<�mҷ�8����9$����h�3�
��5 NS0m�К/�p|�j����ߡ�V�ىA$p���E�!�ɇ�z#��>���q�:�'/.Q�n�\kʃw�p ?n��O��H-x\���`�;�����q�y�B��Y6�q3�9[O�P8oE_A��J���BN�..k��� 3�����%�� 9���r��q��T��|i���Z���O/�ۓ,j	O���KJvUC�yB@����v1d(O���T�8�^T���Οe4����市�,F�QD�A�e黡K*%�N�熱�yd��tG5�Ua3k�(�x;��986�AŤ#��m���
�Tԧ���\:�1(�4p�D�a���x@��Dz#C�Mo�V[�A��
>�;G��#�{���@P�|���^�cOt3;!=�k�"�%�M����i������[� �) �z/�����٨z��d���=�K�#{;jc�������[��O�5qĥ��;��V��T�U�_��Xb�k�<kq]�K�[v�1���D�	�Ya�V���|:���=Hp����[���z�W���GW~�~Ntѳt���j�Jٝtn&�b!�Wv �g�� P'��\b�QzBQ��&�F��-�	몦G�j����18���*���/�FN��K:�rfWrg�
����C�uJZ����^ce��$��h=�1��h�oߥ�:Y�%%�V-i�^b�\��腪�a�ƴ|& ��";6�B5�]-pWd�����"o�O����b��R1j�9�3���i!n�X9PC�M�b�P_tz�`�s�e<T&I�ٔ�� ��x`�=�ڒ���NU��f5�:�yh��:j��%HT��c׆�D�0"��s4n_�%��7�������#���G'��eyg:3J)�6x���{��S�ۊ8ήTK'��
�Ab�xk��S^$ZY &�N>2���=�L�3�Ӛ��.�d{J˙�`�`t�ܻ{�l8���W��	�Ǝ�[dR9��E��33H��X����\l�n��/�_�V��i�Z)Y����{%�_�=N{2w�j��B<�E���+K7	�lz��=�-Ե��_�*Zy��k>=�lqa;,���qpj+�8`�L��'�-f�Q}T��Z�0hx:��1�w�������k�rk��Fw�o�lP^�[`�����#k�<H�V�fq�Ѭ����f� �A�G5�(�mb!�Jq��/�Vb�S֔Č�A�K�58[$�5G�!��7"�f>9�|��y�;r��X/.:Y,8(��4�tA§H�>����2�0�$)��͑t�1&:Z�e�)��,�B�-�%�0|C(3D�c��sVN�T�W�� 	ƥܤF�}�_$�i�^��M5�\�����b)�6�⭈�l�!�����}<��&�i���� զMg��
ӕ�\ ��D0ASDN"IY$��eU�����YR���K�f�������?��	�䆤:����'%�_�����&?I��\�C�3kN�H�Q�>�1-g���ڈ�ʹ����oK�Q(h�2VAR+�4�N���D,o�E��d����#�"7����SF��~iz8M���<[9��ZH�Z
�Bs�ve͚���f��-�牧�D���L��$P��Q�1�I=(ln��c�Iϕ�0�*��'5�8��WU{^�T��ן�v�������]O7JR~�t*`�^��/ͫ�*�$Y���Y���K��gƫ�D���%�5wH�ž�9��P�޳{��;��ܒh3ʱ��oz�/�k���O�zR�?!�(RG֋[?ggV}}I�ׯ�qs�t�!��[�K�0�IR
w�s����s�|���@Z��0�R|)�S��5<�2c�+=l+���(:����	k��W��b���G��ǘ�
 b�<�|�E�3?ܖқ_��3_�g�(צ��ک>��D���		N��~����h
�khO��V����	��xإ%�^�a��~[�y�4�.����b���"$���i���#�[��x��X����������g� F3=��͸�3]�`��.��X�P�#s{۟�����5#6���͛B��R*�Ƽl��͋�������D%�\���V
�N��CA:��!�N_|��%��6ɝ��0Q�OK~3��EQ��1] )c�q�9I�%�VmLH�/��r%���]Z��^��m�M���a��֥
�H�ޏ��.#�����ɣw���y"��̹�Yܤ���6ǡQ��n���s�mi�o$�{~����΁��γ_���V���Go+F�hp~ry��q�����搀O�F�����f�©g���'�3c=�k`E}d%W��8ypS?����m29����^��C+� ��V��S�a#�Y�z�:�#i.�T&ݾbX��/��|Z���}����Q~��i��Imm����#�%)F㎯������)����`�6�5x7X3,S�h�e��2A����m���������-Cv�,{�kY�߼�8��oI�\6���۫Ti�4[�\S\�mRAA�b�Al�U�S$8tfv�:z`��'�N�q���~�(���~�#_�;,���]OkY��\��H�Eo� N���C���v�Dt=I�<�I<Ѣ�:ͷSk?�Kۼ��7��ۑ�@�r!��y!9���S�w�c��|��`���y���Ր�^d�3��ۨW��#�ߣ��|Zf��{븏ly��
XI�%�gzmZ�U�&�d�V̇AE��K��"���AW����bJq�v7��B�S]mu�,��[�/C���C��ad	��
y{���� ��2{�0�������z|퐥;Q\�X�`ēn��L@ܥk#�A�D�^DS8ouV
�M���D�5��C�ˋE�l��uM�p�X��'�(���ϙH���s ��k\G��9��KH��4Y�[}Xw[��������|�ޫ/��L��MkR���� J�ze}�����	��Kq"���s���6c�A[�ţ�j"ܖ�n���ve �Z\Wt�1C�?��X�F�μ)t ������-?W	e�U3$ rGe��u�!���޲$f�͸i/z\���ςB9�Y��M5�23���Z2�&5K����j[�`�/��?��q��,�#����Yws�_IO�����u��b)4�wTqٵ�*�;3I^�/[ǆ������[i���т��xl4(E� 	s���^�T`�{��QS�+�R��}#��l�d�J<4�u����9��t�<T9��/�T}����Fz<��<�Z��=,vl�V��4�舃������F�of�x���g[� ��[�f��?���������P�� �c|��"�~~l��?��B�Y����O��%R�f�o^n�t����4v�?'��h��_��V?c��x�)L; ��*Q�Z���@n�0�P�9�D�$��#�)4����cF�2��{K[+�h�UW=7�g�+A�Հ�7�q\��(���v�����PE,+��>K$(�1�g��vn��n_Ma�lr.u��o�,B����^]S�-����a\xp\�ܵLB�]F�!zŖm[>������J���%,x�m��ùØ=�Yt�V�Dαc<B�  ��E
#/_���Y��Q{!���_uK����$)Z�<�C1S�%����������T9v;��ƃ���({���=|��1����C��0w�0GXJi�|��X�&���\iF�ߪ���4���?�ƺ3�5�P���4D����G����W"r�^|n�v�<qe��| ���L����{���J�e/���@X2�>������z���rVa�������ǃ�r�'^ '}%(�x4ᅬդ�jo��1ėS@�� ��WW��<��>�	��C�� q���xW�.�) 	���̄�����uʻ@���b��o���|�(���E-m����ITrVp㸽��J��jӤ�a�ʖ���ES�>�V�@�u���0��^��$���?��s�ꑨ�)���-̏"BK��n?�nm�/�{
�y���;�Y@y��$�eǟ�A�B��,��:��{��i���*����Lx�jY�8S��n-���O��\�|���f
o-�<�؇h�ߛk���sX��%���
�.�3~��(�w��Hx\S"��&%Nd~��x&"unP�!��֭�hC�x_"-đ'EL�;x�E�W�bcTE���y��3�m��'|ˎ���kbS���!�p����+IF���o��m�V;n��y%����q;�zq((�3��o�|գ�i>${&��1���v�5R�q[����s߃j��0��Uz
W 䦬�%�qI���0 �[<,<�ZK���8�ɑN�q#�#�t������ʎ�d��~����������g�4?�$�N�:t����ϡ.�O����tE�z�2�#��?br`N�	��*������Z��[TЁ�_� z��݌�)5��<	W�ڴћ5�z���d���aYb�B�y,�&�MrE��bB���_^�]���yF˙~�a����˽M��v.��Ӥt���ozWm|�\R��!�`,3a&%i��>��ѐ&"��k���X����X�����?}zo�ˢ�x�@�y�B�l݆��u:�ʼ\M�.�{�T1V���j��%1^��S�Sn97�7�r�:\(4��Z[�/G"�&/4T��ݭQx��v��u����{�5) �Q�X}�E�h�����d`���$|W�yai�a/�_)�� �]��-��"q�Z��9�`���ʖ��5��x�/a��zSP�}��ZگMF|��>*읨G�p��wuh7�"�0�Q��Q�Z�\/]wDC}�����,a ��E4";�.���b������05@=*�XG�{�<�
�>u�(��������	7!����t]{	��[R&�o~�N�#��r�,�J#tm�����m���	g��m����lfέ�2Y��0�`W�cE��緃��F|PR�(���l$�t���f�[��G�iޫ�U	��j_nl��5}�}�T^g��)@zݓ��4h�"_����.��׬-Vɪ�v8��4.��\�ϜN7 ̵���qO���$\(��mg�}&��m�#Rv��r�������ĭPn�3֊#gR� P�Z� @�P<�C���9�߃����/�.���`���,���vR�?��e���;9u�K�z1sm����]���rXU�H���'av�	�� t{�p��}׮u�e�j�&�����^N!m��8W�KdY��������5���Q�����jJ���M�-w��]2nt��#	?���b^��W�!�+K�/��@'�w��M��C�E�/S[�m�@���(U;IhE2�h+>R����cK!;1@A ��Q9�W5� ��X8�7	O	��z�Q�B�	^}9����Y��v�x��J����j��mI;�`" ��r8H-��5x1��{" ��Y8���Qm�A�Q1�K0�$9�>?6����7*1T{���x�� �_	I��)*� "2�=�@��;:`C����?���|��͎�ڞ;SW 5b:��y�:	�QCW�T�k�&$.NIw	{�u��hv�"��qe��f1�CPh�߫���y׎���������6��g�,��|�P�m�<P���X��|�O��(W���ax�`�N�ޙ�Pp�q�݁xXI��2�b��	X^�%/]\ӟ9q Wb�Ip�2���m�82�Z�֛|�=�ڤ�lhx�X*����Ej{���ºI����@�n�D��!�*�7�@�45�o�{(�М�T��o��hP���@���/���:��r��S�px��[����|�1��T�7���?��?=��M����]޳dq�B�L����$�*4�
1��Ŀ��p�u�
���Q�t���Í%:A��� Rs`Άbl֥|�GN2n��d=_��ԡ�ڧ�~fW�r�X���1'm�S�V�5j��B�ܛ�r6��L����fܑ6m���
V�2ԩU|Fø�'�E<6C*♼j�</��D+�>��9iF���o-�'�xi��s�#ݘJ��]�a�B$q��e���ٻb/5���v����7Lu~�<iY�(��s�J��
�Be��mz"\���B�Ma���Qv��UJr@�U�5ObR�!���_)��=��}:a�	OIp&���.�3r��=h�
�R���^���nd��r��h2��C
Wh����b��I��h��#�N��Zɐ}�<�lͬLw����F����PG��e�p�vzF�u\�5�6��
V"��)����t�Q�1�Bm]:u%��XF��rYG��Vkt��+<����I�uv;<���)w��D�qQ��� ���.l8�h1��i?E���o����=h���u����?�7��NAU�9�>'��YAY��y�w���,;�ϳnCY!�����û+�R8��a��`�ž��P8:N$�_�Ԯ���V�) A'+�G,b���Y�Tp�Ϡ����{a�1K?�?�t� �7�僼�t��+������<a���6��u���M�}	��.�d�E��0Fa����/��ӭI�P7��d;I���g�?܇@�&F�u�D,�@튭~B�]L)�}׭���?����wU9����h��
�Z��e�:]��5m�w�Y�V�����;�H�(�_��+�0��&�it�M�I+|`K�T��Z�Q[��� @O�GT�5Z�n�G99 B7��v�s�U���m�3�{���r(�go\��h2=0���wh��=�;���2�*S O�%M,z�h�i*��W�}���da0+*����N�'.P�̈lU�����tb�+�P̰��HW�Uz��Z<$�)�] �<���jR(�l��:}\{	#`��$n`o*]N�l��|;�P6�6r�&����}�Q~p�:v�y����<���n���$M)~ ��a�AbE)�.��($Ѧ]��(�En}�	 `�q���&������f�3uǀ8!%�}E���0��$jR����v��6�Tx���M�@U	��M��V�@̭��cO@�4�u���|ӹ��ץ-$�2����������Vj���3y�P��s�r'���(v�4��i*s�v�e�J>�N�>��([�*��p��P\ۏ��݅vԶf��P�Zd����U�L� 0^��m>�w5/&3����5�2��<#��3萘 �uB>�����7���MKK�e���N�J���O��7a{� �z�(aU�,��kH$K8��]��J��<��׊�q�9�7]*�f�D7gG�[�MU_=�%� z�GUѫ�^��X�	L:��y����H�Ԅ���胦5�rt�O��Q���{U������ڹi;)�gv*(jV��0����pn�{�g��[$i��}�yRT٪L�{O?*�dVp��1�D������%�(�1�����kb�;�]���"[a�|*^\�R�=պ�O��a�Bk�MQ��5=g�
��d���uH�i
=���Ys��:?�,�=g��M�<6W����e+�k�"5r?A�����c�.��~val��x��������#��]���C�@A��f�	^p���@�_'�Y{�AS%�O��R܏D����7�0���dOġ�|/>P#W��(ȃ��\*���_K��Ka�
}��O%�bv~o�3�2�?� '��zZ���Wڎ�%2�^����o�`�ȵ���L7�c߈C�e]4"h�-Q�[IC*뭥k���s20��Bd�㱥�;�p)H�!��WU���RLe�T� �I>������㹏�����\����/��NT�uQ,�`E�uB?��n�'	�&��D�!����@Np��GFp3:ZC�X��rqyq�6�mK���%�k��ŘP2���r�O�-!7õA�يKD49n�O]�Ch�P�x}���9+��?�p���s��Y/�������2H����H2�ž�A��N����_mn��tC깺���TӨчq>�e]�8p��=т�6��ʣ�k����tǦ�g��Sr%q2��TC�Uy�,�5:�� �I�Ϩ<43~�.7�p&�.���Ǩ1�I��#T&>�o����lg�1/k&�< �T�xn�֏�
�l�1u�fY-͊U@� .��{��(j��>1V��f�UOf�Sq	�iRd������#��h�o�j��A>�/��΋���)�?�1�(F�o��I�0�8
���(�p�8JiL@Z�Jo�0^q@�2����{	�����&X�ȺB�b�i-����zo#}��bv�t��O�!G�~16�v	�pت��5XU�e�z��k��pOqaβ���ʰ�і�q����L�ģ�C�r�{m(/f�^@�S�� ��<1a���^�+9�#7dPv�7q(����A�[C�RL��{o�Lj[��E4�"��I��&���[�~х,K)����L5G����{Y�{n�H����]=�c�~̑д�co�މBg#]�N��C�@ӻ;�-�T�$4e�����J��"!�?
A���\8bKv$#�d�I˥�[�[��k�Q_����}�Vy����&�����(T�/`}8�B�e�3�Aq]���MKe�����1	VX'G|Γ����Uaڧ􃤨�������w�>7+�)4��dV����=c���,u�/k缌�=���_�$+�$�" -1+��$�Q�D<�5��4H�a]�Ӗ��4�=!
�b��A��5��[���y��`)T�YS��4O	�u����R'�m�̥�m����aK1A�P�_�{����[�c��Dcx��L�υ�T<���rf�X@�}���7d�N ��u_|"��?�}0z`���==�P������<�?A[����é(9������h
��ĵ�w1�R_�0�M�g����f����\��μ->�o yoŗ_��U�B%m�y)4� :� �}�����W�k�1%��V<f��n��n��2&b�����D�%biN��%��]|U����6�L�R��ޡ�!u.�����ԆJ��H@��O��6�r�;w�ЧͷA���|�-6'�j+�"u0��ļ��~ҶZ6����K4m��=o �2ʅ�]GJ��:���kL�_��.6�u0HR"^����Mh=[��W�h�� "@�%��>��O 2ƫf�j�_Zõj��2T��c��Z"~�&.j���]����l����o����O(	~Iֻf���'$�HC�4-[�<槖��2�_���%��̀�U~^E���:*��ͭ��o-�jɸ�"��4�t�5]G�Y�)k�]�'�r�	 h�|&��Ţ�m�(�h���x,�?܂�����5�1�q�7��\[�}������Ե�v��r?�ݩ�0�P�B�$���>��v�-l����f4U��.Y�F�>���c%�2;�5�9�C[��:��'MS�J�;���g����`K]Ӱjxtl�OE���lP��>��2&���S�;�ާ�7�i����g��KZ:0�(~@�+_��#r���^:ޟT ������RA��<�-9��x��+�\�`Q� ���ބ0d�/��KΐWV��4t�Cz�<lۀ�jShP=�I-�J`Q���X�$�\׳�'q���B�&8Qj=�����~4��6��\�H�k��� ��}�����}wF6�u	�d=���L�K�׻H� �JcTμ�MϢd��[�%bxR)'�~"c�
}�:J��(��T�N~8%�����,���%�s�J=��~BlĪ�'��~alA�����.sw-�Nt�������"�[�4���O�Z
�y˯
m�*Ol��s��.�0e����x����2w���e(Q�9�5?�=tD��y��̸�9RU7���T{�l��a����b�U��Ē�97�A��Ma<���X)����x����H,l/��0:��(��T%>n��|7�
5���qE����cd��^"�w �Q�����aK�>�bY��j�"8�0�R	�{�׺{�eo��
?x��H�.P����`}XS#V�k����c/F�%�� :?IIU�I���㿕��ƕ�R��W��P؞�J���F����P����۪U�\N��&�����u���e삄�M���qm=!������n�Š��x��֠p)8ߗ�w��A
	0o�,�~h����4��Z���|ʪh]e���o�]�)���_ӟ��:�D��� ��Ɋ5�n���VO\8�
�����\�n�cҢRZoej��b6As���H���n!��B��t�	 <�%�0���D�BO���<oq�n<S�/��{�p����p}��W���a� �H�������N��K�]'�@6�B��6�+�)N�uȯ:>A����#ؠà�A����iW��ҙ�����XD��'�:�W+�w�G�@���~��P�]�h�T'7����#�1/����X���� �"���O��r2��f]F�\DO0g!���/b���o�_��M�;�T'�z�2gb
�_���n/an5��)�w<��ts|BK�5hY�`�����p��=�/��6�B����|)ҩ��na�fJمQ؍6ݐ'W<4����"�juJP��SK�|X������L�N���O�� 3��T�a0r`����j����r7'�-k�J6ziw2�_�*�x�X���z��=�[��	XR���gJn��CFG��><���Y�xSz��I����A�F"$�����^@��MS.�F}5�.4�YH��?:&�0��Z�7f�pW.�����Љu����Y��u8���0:�鹹ȫ�&/�PYy.m"W��H��nQ{#c�廳n�*^�/��8�HM�CW����xW���enp����b���
h���x�
E�$���PӮ�������+.�1�&�1�qۤ,4�	{(�Ω�G� �}�6�mL~�'�9_1 �}��כ�n��i�U��/�M����$* (��J�1���U�,�ta�uDh�����R�����nG^���hsT��th���6��D�6���<*&#ߑe-s5�xIE���N͋����V���P�_HT2!��2��8�K��E��,{�Ws'�n'�.PX�| �O{�]D�<�A�'r(y�HC�c��){χ����1�-�#o~�'h72m��S�V=i���x��g�C�\$��T�[}cq-hy]ؿ�&Qm��ʠ��Q.|�����i�U;��B:�>����- ب��.�ٱ�4 �� Nh�N�I��N��!�S���𴢷�%+d��?��y	�!���D0�0�|��>ȩUg0�m-M!��n���\91C.k���شj���>�x��,�pI�I/�p�	����8�Y31R�,� �]T���Y3�($ɹ�k%J9�J=�آ@Nj=格L���l�iB�ీ0�� �Lwm|��sM(��3F���v�8j�:���~���z_{z�f�]�oi%\��hWy�$! D��n[OQS�.�5���3�r1`���Pj�Wn��X@��SM<�X�G�T�^#�_m�m�V	�4������[�OݼI���Z��m��l��b�59���]e�-�jXEI!��Q���l��˾˸g��\Cʜĭ]�.)�4R@g��:��.�]t� d-N���7�j��}ֳu�f$A��� �>m;�V�ݺ��I���ڀ��Fr�
�%q?m���/�o��+�	��O|�� %p���M����ӎ����dIo��$��*��>�W��[�|�ԍ�����1(�n��,�=��e�_�yb��ݵ�ɬ�e|�~G\�=��ZÐ�zʾ�	1��nAQe$�x]��
�pq��HU���F�h?�!��	��d��*띚v�/���Z�s�y�;<X��*d�`�F��Nޱ�Y��.V�4�ͫF�bÛC�|�B<c�+��n�מ���8�G_�D�g�h��]�n�B���V�B(_J�ͺ��F*e�^ɱ%�[=��b�%4r���&$Ȣ�7v�~�]{��kغ=8�b�H&�Y��Ra>�ܩ�f�Uǒ�x���.=`06�b�n�sr�&�6�3f2��C֬@�+��R��&H?��j�����Ī5���������߆�z��M����n�I]Be��a|�X�0ŗ��3x,  Ӌ&&v�{��Pr������''+��R'd�@q�����c�,�	﾿*�,vւ��(
m��ry��XyvwKO&iU,L��< lG]�v/���g�'����k�]#i	ř�FWl����c�kC��P�����L �䨨���{��H��nڈ+�(�1���*3e���rL=j�Dc���كMF�~d��<X�J���̢+�Jħ��l�a��>��e )�0��X쐹oS�6�b�\%�����r����w�>A���KE�\z���傟��zI���'���wf1t�����W������Ŋ>��ʝg`�47�A��[1U^��A��u6��cH�Z�i*��>q�G�ϐ?��ٵ$(��#�6��2���?aU�C�d��s�8=_�. 6=D�b�4�Kv�}����&ѷ��\��Y��u ���_hk��9��#81�[b��l��86HIS��G�����jח���!��46��H��'��}���^X������Ť�R�=|��D!�> =��I�t������/�&�q9�Y
��tˆyx�`���?Oz��k�c�FM�G�	�:m�w�+%�m���5ic���Č��_x?밵cYxd����9�o�zF��A�И}Uܝ�G���bWy��x�mĖdp��0R�p�X�p��XA_JFtc�7�����Q��/�n��2O��C���pY��y�������O��qO�P"��I*���>�s�X"����V�e;9�H����Zd� ���\�y}�FфE֔�����npv<h�d�/���V��q��|9T�����.^a]�I��Β�S=��(���nf��׹A��hz6�̶q��om���Ô��!�ѵ�v�|���$��|��n�HS?��FH5ٳ%fa����u�$VoQY(���f�i��r����o�?���x\���#$�4-��\{Rg���b)���.gS� ��f6�4�\D4'���r�Lm,c֎�����Q 5M�=
�V	��*ԯ���E2fX�������W@�KdǗ"}��^��z����¥����?@욛�8aU{����f�L��G6���q��N+.�b� � .�Q�\v�5�]�o��\e�0�ǹ9E@`��X¸0�.�yG��rʒ��B����e���!@{?��?y�v�;s�YM-G�L����G�zw
x	���S�&�`���É��y;��8H-���B��)�p��ǋF_%�U���l�<-�����e�ƁK�A��w8���=�L2G��sR���(�j8�+�wm�5�r��?
' ��<LX'{B_�<~�vz!0�_�+r"�U�x� +��I\˯��[_)�}�s�y�U�+-U�����n��5�EVE�`n�I�̫�P��?�e���q�,���j��mRI?$����Xe__ԁL�g_Q�.�y����,5^�0��tl���_:T/&Т�m[�p/�MKw6S\���]�*�� T!.��;���a�[�������傩�y�D�qXIɈ*��S��\�Lpj-��	v�.]�݆ v�b���^@��8��1���@*�7���켏����<_Ҏ����l-#�7�S	�P�T'R������Y�+���*y�`֟�N7^�1�6D0A@��)��5�ܮ��.L:u�R�q���u�`�X�3>�>��֌�Հ�/�w|������@��izHj�@�1x�I�Uk�b,����w��K�w���E�_��.�K�d}J�~��
�#!!���X4��g�P��FvJ`B����m�vZ����#!��Ix�-y=9��P�p����m�Nm=>��Y9�|��(C޿��K�Ȩ5�2�{��`S��.�4s�3�yɤ�A���凧/���4O����DD:P=��v�0x��<ك.3Ԋ��Ud�~\wx^�gb�H�7+��]�����18=6�d�E���V��:�Xao|�������\(h��_2L�+\}�5޲*��'��~���7\t2�o���ib��XQB"�b�_v�����|�M�D��	.��&�CHˮ�o�ո����v�eI��|T�ʹKuV�P��oO��!�-5���&gr0d�N��7��:��G��ڨK�,���4Z�(2_�^���������x�א1s��DB	j����P?����������
}�v��P��ϐ򟩎��s��N�lm7<���K�!�JR���xg�*���[p��Z{�F��X �'7�3d����� <s�8�<���m:@��ĩ>��<�LK�֊�ՠȉ�l��N!�F1�ݟ��!��IW�[�j��Bp1���U��^
ɞ��[���ɔ)fú��>���)M�o�/wW`L��B�wޤ&�/�ق�qL�����(�.Ñb�(+�W�>�r��N�EHB�y�:�:��KZ�q����pp�<��v����L�N�>�2SY*��K偣�F%k��G�p�M�!���Ӷ�̗Z'|E`gU��_��z�#�Js;���	v��v-l�U\������a���j������y��扺m�48�%6m�S�ih�D��GtTe���b���|�́H��Ü�f3�.�d�`U�a.
�T��R[��(��)s�&�	�R)]�@2��c���iW��	]}ӛG��9*P�ؑXPk}��(�!9��m���M�
����G�#3�v���V��d�2�/S����>��1���7��� /��Y��B�O �NxFa��h�];�b�
3��s���$
�)��rZu��so��澌��Mi�5 � O^^��!U5������b��WE"aO?]¤�<m�	�O��q_C�G�h��
Zzb>��b"�3�X�|�G�6��� #k0�h�x�m��_��	e�ԡ^�BiXLqgY;H���vj7y=���zgѲ��N�=5p���3����+4��h#���z�h����ysٔfҒ�u����&GA�	 ��Q!'2�u+�E%�F�E�I6��7i�h�E	���`�>	�n���ɫq>�V�qpdɠ��g`�gM�#8��c����-�2(5��n��>��R�qa���oY����k����Ŕj�,{�v�=��ڣ.��F]���`o�=�\�8a��]����=����x���4K	2F�Q闳 OI��8�16l
�$tj��`H�m:b�dծ �'S-s<&IrA�-3QY�^���!�z�c~r��5|��|�)uQ�@>v�B�\�0x�������"\=�b��7̵���فNo�~� ź�ޠI�X{O�r��N�~�u�g��� ���y"f^G<#��_p:��Q��ס��lV����n1.��ƺbԂ��xD��fV�HB\����JY�V9c7&��NO߭T��Ʊ��j�^`j�����:0;��$w���ë� �W�l��b)��7B���&`�:\qWv�0��B]�L�
��49ވA<T@"�b�>4
����J�'����c��:`*�#z{��ԏ}w*D�,��H���v[˳ ~ӕ��	(�m�4u>A��'㗬��W+��L��}���|���~�n�����jr���Q~(�$�#�I~�����L�O����]�F���&��H�,G�������e����6m�ND+n�į��W��W������'z5�aO�K��_g<Wſ�(t�6z%�|Zv9Ǚt
�Y�ϝ���,d�i����mR�[7&}�-��U=GǇ�b���o����I��3�?�ߧA�/���I��q�V�8|�4i�_�^O�b��;d���u��|w�(���4���@Q�
��k�3ˍ�-B�3@��NC@�	�r׸� *}�\~h�olc���;'s߯鄏��v���R�&j��(�'��<:U��?�Ǣ���=`
���k��%��!h���]A)�P�*ݾ�.;����'j���މy���2 �,a�hbȌ��@e��цZ�r��R�l�+/���eq4c6���ᰇ%�L�� .���;�!~82� o
6$�Q�7�4��Ҁ6PDtY��DMG�� �*$��	�(���31*j�X��I�A�����j��3�	�QG�j���P�5��9#���Tf3g�Ƹ�,��Z�!�~�=1���1���a�-yU��]�i֢�	7>,�*a)L����oZ�E�{�,q�`~)��LevM[�s�"��ħ�Pn6@[E��'n3�v<�J	#t\ˊ5y�K]V��G�<��"]��4?���,�8)�-�wח*e�MU��Yb�&ܗ��N��\��Hnԝ/[i��i�����W�2�x��:9 m[I��)c2���;in^��-u"D��N�8��e��=}`�)�U~j�8 ���b��>������e�a�|�!�-�g4dnT���ۛr�I�gc�ky�V�v��@�@G�u?u�Z?Ե}n��2bz�JTv�&��#�}i��'�XV��Fh���~��Ⱦ0��^��	A�,{Iݳ��XG/�@{:�fP�����Tl��w��CQ��{+�q�uR�N��v��'o�^"b��6�|r�Тf��Χ�'УHI�#�QK�}�y��5qo�|�l���Y����"
��=7�'H��}�Re8�u��>8�����s����<�_�J�6�K�7���z?�^��^f ��iS�@VO$&�
���h/� �v��見���f�8�M���I%�a<����3��	$��`f/]F}�9�JRs�(��$v�wܕ;���mX��w��r��j�z��Cnz�XO�d�������u��_�ٹk�* }?֭r�lf�o'�Xŝe)�%�_4�������(�#}'�.�Wx|��6}"�$�69fF����wd�MQT'X�C{%�USR=����ݗy��\8NT"ؿ�=��A?-�S�X��6l����duŔ��XN�Ğ�(oB�
x�󌢃��$h\߿=O���� gcߞ2ê �eT�8<�;��_���2$%�~bܬ���V���I)e��B�Dq����.z>�!w�L�L��]��	ZE�v�D0Q�0<F��=���I�[�~�j�ir�<�.��70�g��޼xF���Č����ѽ_��x����&�NX�ߤ���9O"7:y������z�:)�F[��]��"���^4^��l������Q��t�V�!T
Ѳ_d�2O�<̖QJvV}M��<3�j�o<o����U�&=3��|	���+�8���u�/�|N����>�t���o����*b�JSE����P��1f4��w�t�P����pjN�?Re�xM�J���U��J�i��Oft�	vm��I�ܺ�"���f�?\:�a��=a�V�!�A�'�e�% f9�>��Q�1^�=VT&p�D�%�k|��aqMׇ��gY�aO`�bGfxi�u~JPʃ(	L�&Q~oC{��s;�<#�j�����8���vz�H(��IrL�����l��x6�T2ˤ��iok4 .S�>r��@�ʘ�Wk|7=�c���W	k��J҇�.y�<8{���K}���Z��f��Թ���&�W��U�y�:��t��	�L�ē+6�-���,�-�{�b!�.���!̓��w僇�pW�ǽj=x�
��=O�����eJ�;���;����U�G�dY(�M4�&�8���)2�C�xE�_1M]��&y��c�ٙ�؊��9]�j���(����D��pX�K���m�;�o���
>�%/��""`��O����ù�zG�a��8,-ŵg�{��W���nK(��}��������".I�}�{r�!���Mo=��_D!I�\^�*�}�]��;��&�V/��=b:."e�1(�yo��!*�����d�_�:(`��7��dݧ_;�W�&�ډ�i��K�gx�ԋ@��0CBFL��� S�(�M'7��Y���cRz
Y�8Q�\��u0=)��T%AW.�|����q�¦f�^���<Y	N��ښ/��Ib.��z��~^&k�g˲�����T��ƒ�����;O����@@r=BV�;7~W�Ke���r���x�r�@�%��w״Iݣ���!�K�4j9'�q>l�F��,x�~�ٮl���
Yuq6�?��]����(���Ǵ(c,>D=�oۇ�ae��k5͙�&6���ۜ�C�fo_r��%W�׈�(��Z���}�ݞC�)����Ϝ����٧�-+u(P��$����㟯��#(��������}���8=���|��V�6��֌K�E�d���R�ȏ/!�]�f��#���1�)����nd������/G.���M��E����G�
�#	�&�����f�׿MT�,L���*q"VOw���wrs�Y��q� -9��p�FZ{�m��\ɭ��|<ndb�� �)�u�/�k}�7�BH��c���qL�k��O�+���XjK�<��1� ������Ě]��$��j��+��J2�֜�)�\�o�:���̴�W���T��o|��X��K3͓�y�kD���F$ ;"eԻ�����)��G3
���~0�W�[�>�ܙ���|������8�>��O�"dr�>���ҷm[���D���#��[�����&�`@3f=�%^9'��F)���};��\de�zC�^��� ~�m6���v�BŚ�:=A�z�A��@=�������,�GOf�Fi�n�d^�+������O}`r���x˼��Qoe�.EwX#��,Ι��"%���4��t��hm3Ě�`d�:Pyn�"jo��Jc��BР7'��E�Y~��H�ׯ�1o�z�Y7H��#�j
���{)�tg6'/Tp2|g��rPF�f&6�1r��?�'S��^��vB���#�n�F�s�����O�Q��`ݻ=,��e����\1�!Qb�EN��i�R}�b5�;���;��^�W��ڸ~�9�	ط|7�2_D���g�?�9b���*5���TVɌQ���8�f�V/!�`.�~^�=�	���R��9Gg��p#_�c��M"B�/�闥E���T�˖�������7�d��׌�l:	����cH�E�&l�*[�o��V2�i�	/������BƲ*<!��ܞO��m�/�-��H�l����ʿG��K�O\F 
�,�P�Xf�����I��=7G/�� ��N��������>J�2!��cd3J�IieA(/CM©@FYH�y)��ĄtqP(W�\���`�L����EC�őddH45U���L�e!���P��=��
�x6nӳ��b��������P���|/݂��e�	伙xu���S��T-�(�n^����4���y\_:� @TOk�\����O~ެv[#Eeͣ٠���cz����%�N��TF�&��n�����/G���F�Y/�S�LB#�kt:�u�["�L����e���J%�;s���p �ĺd|kn�uTmY�W�'����r)y]���+�ˇ��F�B��i2�0��*��n����
�xo]�k�l�GxW�JUYƴ?�4U_ �uP�[�}�#�A�NA���h<��R� 7 �l���&�������8Q�_ԣp�ik�X2�S�@��Q� �� ]^�F���g��@�n��?gQ�5ߚ�#D誝��_;-Y�����P�����A���ӛ5�~[K�.QB~�:��>����f��q`ʹ6���/�{l�"��˱/�H�I��:�_?ƺ%�!����T$���A�c��j�G����$����ka@���9���"�E��K����p�h���,�K�9���s~N�<�����L@]�a�òb��&^���b��Uo�^�t�GsN�'���;�u�#�i	Z��h��c���F��b�鸹�����}��O��<������{%� �Fi֦�|Z;��oM-�Ũ�(�<N�q'�z�	�k�١� ����x�����p &#W9�OD�{��� �g�n���Ѕ{��FX%��ߕ\C��_t*�rEl��:J�*��
�,��e�w������������`o�@�������\����ޙR9+�<������U�
����D�o��'%�G�����q�e�v\ד� h�֑�\�3H�u����CQl\��a�o�e6�^������؂��75]YR�~���+�#�k�툣(�֊ ��in�_�����5�o��>Ƭ��s�} ��.q��j��@[Ħ�/7�XF{嶺M#��t�G��
,T]f#�.b���{-Ycb�=��S&�U��@M��^	���Ӯ6mi,��W@�%�LZv*P⏖��w�P�����Q��3X�4��$�����ޚ���)`���"��͊�N;Ő�:�P�dL]6VYf�N��e#�����*IU|t�ꟑh�P$���9�94��1>UĄr�!�4�u`�xN��VX�}�f��(l�&��Q�Y��s��%���yf⪟t���q��>8?�;�x��We/���Kn���]��2ضWH�!��*vrq��ԙշ}�H�y`!�V!��%1�_�{Y�mO��
�Zy, u��`�L�R�B��N]����Ꝉ�-n.��` �kG=zG��-��{�y���蔚ߩX�|�2�k̥��ʓk�wpR>y�d��4*�^�o1&�\��86�xY��AΞ���v��,��^h�v�y��V����~�w�E+J��~T�=I';V'�B������b��_����>�1�`#�	�/}K<D�Y��̀�ds�~�L������Fi017g�7�� ���4��3��ߙ�^�.C�2��_ѹ2���a%_��<I��������:}�>���Oey�j�-��\����|އ�}�+i�_�?�꛱����}���d�3py���ᘾ��+F�6�[>ϓ$!psg�8:?��������$*��-^�#?~�Nf��y�u6_���7�\G�Z >@�ֺi��`�#�a�O᪟Z�>��Y�_�n��G��!��D��7o�ܽ�D�Nb�}�\�e=�Q��J�i��V���}Cd��ڷH�[^�붘��Ţŧ�0�Qem|i)�$�a��D� p����O; P�l��jC�co 	h�0����3�/�����L���KF�!)k��ns�����Kkae&�>���k��?+C�ܥ=�#����Oc6*�\�ֻL{�G��9ݟ�8����y�?{H�Z�$O��0�R����,^`UǛ\< ��?�`.)�A�O{<�BϺ��GC�.!�t
cU����1\��S�3�b��	��v�Ob��*��a�^�#?����\�H��O�����D\>��s;Xԩ�6��� ����uC䜚[�9�T�Q-���q��a>����B���>���/x�4K$�����󨉻�_8�}���,+n���Ȝ�
BI	e��4�d3�P�������V���GM�ɉ�N��^!�F��s�<�טp7�!�ĺ�%�7�b�k�@�Ň]�p��3�zt����@�e���g��|���/<�P��Ԑ��������"��q;��f'�\y�̼�g0�)>�ʓ�-g�c�C�I�<3��"Ii逴UI,�Z�=O��I�����:��0�OUø6��5�_������K����)�(��7�HS���u�^ѫ�N� �9&YrK����,��_�"��*�7'�J�r��z���k��h��i<Pң�h"Bq#+!��e��Y�f��s����Y8�<�	^B
����k����-�A1XL6�%�NC���լ��HOBwf���,lӰ����ZjS���I� I�����D�au�V�ktPn�eedș}$�� +�ت]I�"p�?X��dx�*�s�9u[�j�\F����z	����4����z�B��wߎoWI.�gm��d�#Y�>c���)��>�����^iOK�/ccI��8�e�s
�Qn2*̓P�q���;	p�3�"o}�z�
��f@��hQ{�0 ���^�'��M�e�/T�yKuP�k�xÿxP5��_��WP�?���%� iVwq+.X�]��J�k�1ϺC��
��z��~�����RI�g���&�c�<���w��6)�yQ*/���`Z�����8r���\*U���?��X;L��ʐ*�qQej�S�WO[��񳴠��'����b�^YVٸ{��U����Ŵ�>���Ϳ�l���@��0Gt�~,�C�\�̃f-�����x������������Iv�?����}��j �9\�ke���.��4�.��Qz+�sluѫs� -�|ݾ=�s�ڲ[RLk�=��+�n��6G��������G�xR��C����o2�@���`��T���y��� 2F��wl����h?ף�?�ҕ�� ��b����
������'6�4�[�,�����K�O��l��uvA���5��&������= prE���4��~Q�b[@�7I�7,���[���)�Rm�,��.$3X�ur�AXA����!���I��k���D�D#*�dp�d��2x@Cվ�p�f��9��,���۸��L�q�Z�u��v/�t.�1����&�q]��Z1oҾEG�g�_��*���z�:����TG�V|�f�ʑ����9�V4�dҝ�?�\��A=��{�\	dK���Mٗ��Rf���#�����ynV�fQT�u5��	��R5�`lS��x<�xڽ$�F\�ѐ�Z�@<m�����%t}��IJN�V$��i'j6�;�N�Ⲿi�6��4���c�I|��p>�Q��WSxړf�rI�l�p�2шXݒ���������bx:mM��%��M�"��)���R��CE��s�4'�I�E$�����^#�U΀�w�\����b��X��TXM��b��A$��62e�<!i�ԁ㜍��	�0ɣ��%��m��������j�7��y�ޮ�;d։;��Z���bO
Ē"��}`d�u"��_�O
�`b����@�ʑ�!�S���(�o�X|�{�O"��4sS�8z�*�ZbZ:^l�ߐ���z���4]H^O�����+)K9C���{߻!}ilA�&�q� ��'�d���u{�B�S���?,�)�o,xM7�L2�g�TH&C�yQoyP�I��^�)�N1pQF���G?w4��u��wg��W��<�'�fc��]�d����4���4]J�r���<�x3O<�b�"*�!��زCI峖T�G��s�G[֖M�Qn�rr�(+�CO���LC�ys��;'3D`����Q��i��0��m*�ئ��f���;�p�w�A�isf?�1���\;-��A>c��]hB������As�䥊RE��n6$��sv����4ũ��-*xb���$�(�ϋ� %s�*�?�Q�����ü�x�|�M�ǡ���r�mw�����E�vI�2��ˣù�H���H��3,��5�w;�{�n���Fq���q��6!󎻽l�m�b{���i�b�ӎ���B�|���[�E�rr�'Q�����ſg"�Hͳ�8��+��#i�5x�O|�l�]�l�X�ڨ���g� �; DY�4Zg�~M@��O��z�|h�@*��]I��ʬS��h`~商���E��B��XM���Kn��׋��ġŹzh��ٳй��e�覨�A�����[w�,�� �e(��ˠ%��[ҹ���d���^���~�v�7W|���y�#I���}&��V|w�|f���6��6�.���l�*1�T�v��nLb��pN�|6{�!�6@�ȏ72���~Vs����n�
�ߩq�^�T(��쿇U�J�5�0f��&OX����:�%�B����sj;s/�%�*Q������I��W��L�ٶ���}�)��D<d=Q�������T7P�g��W{�uY(�m�.g�l��
��d�^C�W\x�ذ�e����ml�H��j_}J�uU�ЈРѕ��n�������ӓ�'�g���t�)�UNH|��rS	)��l�}��Ѓ��*q�V��_�#�6�u�Z���P`�;����͋$��ձ�<ނv3�v�o[o_�TY������H$��T0�w��~ju�0��?N�7tU����h.R�p��0觀�Jio.��*�-3�nqF{�$����'�6�j��a��p$��9������ĕ�0��V!r�(n�����Cģ�^�� V��+�؃cT�3"����`���o�P$Y�񲤂�\�h�<~���f��H���-�}f�!�ʉ��2=�e��7<F�1S�<fJ��nx���^7�rY8<����b}��a��\���m�	Ë7�g����� �9�����>�28�ftNb�to���,�pw��xj��sᇩ��u��N�IK��Wy���31��n-F�|3�N̾�L����cȓ[*�~|���QF�i��Pj$84�7#]���q��tH�x��h	1|+?��tK���}[P/��-��^C�i�+�\�oXK����0�g�(�%;Lc�Rۖ��T�� ����(����B�qŻ��1އ.���{6m��3�����\/�	eee�/k�F��fT.v\����%�dUvK�X����.=�� 9��TarFo��l�^��֔v���3�VR=�Mt)Hyu�ҍ��F�8��y{l���Q���ꌜ�32��qh�DW�Xb$���C�;Ծ?��2��ۋJ\����P�ռb���,u�7[NÌ��6�0g��ƌ�U�g-F*._&Qپ���������z��78�1-��- 3��ݰZ;Z_���������������1ɋ�a|*oY'��7�Uu;y�֠�i]Jh�z<���X� %k�ӍF�E��a���\�����i�Ӊ�s�}_�q�R���<�%����V2j�0G�2#䚁�
�O���v�r�Mg�e�� �VEK�����Q�F�yޒ��+����ս�L�4P����6+�xsvZ卣�B�����򓠵B��tf��hs�x���KK�J�J=r,� �7�������W��jP����y!^ɍ_e%��Zu+�I\^J	s���F�	-��DS��R�!�)�r����W��.��rK�� V���g��V o��F G�Un��]��:E�چ�&�n��Xp���ZV�T��F�I\ T��z~;��]ؒ0>�Z�^q��Q����,�߽�;t�j�v���?L�+l�ܜe �4�~9nA��V��_�Tw���R�1��S/[��k����g�+�!J�ىt��Ʋi
���8/�L~"�<�Щ��S�sd����d��׊�g�kD�`ip��k��K�޶���]m� ��J�f�t^����Q3���ː��=^�<%�����{�
��Oa�O6��1Ծ����ު�/�5�����x�g��)�~�X�s�0%ai� m��٭(.��Ts�^��9�+1��P�A�O��I9�!�����t�7�.	Чv�����m{�=�mN �0����h���؇T�aF⎸��_�1��u��q}<��J�y�z�#۸K�{����bC��Jz��xs/��Ԯ��sQ1���=n\܃�(p�/�s/���'K]�����,�v���#����i���F�F(1�o��U��%��_1>d��1x����Dl&�4���ipduT���/ڏa��Lk��`?&��^��3��n('���Ɣ��'����,No~�ݑRi��b�^��ZBդ�2sm��-�,��pe������/�C^׈DI�h�pp��G���|��w���d�;��.��"�^�,�K!�~c�%�2ԧ�BR:�i�:ŝE ����~3�Y��g}�d��S���^Wu��_�/`j�~b���R�֒]M�?�j�J�0S�޸H�V�r��b�v�U���t�͜�\�X�Ib*$��7g���kk�'?ڐ�Z�m7FU���C���sJ�:�k��4qz�;M H��YUY3����^q|@]�iJXp�sw7nl��e�1��d �J��!S_G"�w>>t���Y�NFr�7�HM� t-��������L$8�h�K\�����UL*�》BI�hY�"f�D���6���ԓ9����,��pYr��,�}�\�Q&���/���s��3U��}�#�@v�\��(��&�n���s�A�x< )�xm;�9�p��u+h�ͪXh�$r,9��_�	�j�eh��zN�d���qdl���K������Cק�L?>�gƈ���,�49��K���;�� �ЭL�L- 2��9	��cj)��e�\F���i5p��x�!��������.��9�ð��sg��k
�?@�j��[�=�4R/>����"��m܆��<��A���sb-�	�׾�\�G��9�B���ɀA�r��fSx'��K��_�D1\�g�Z��ȶߪW�|�~�ܓJl�MVk�GY��B���^$hӍq�ɒ�w�p�n�e�9?����X��еt%�:+�b��^�}��.�eq1[�Ht�+!2�#�6���N���D2T�]��
mMNy�6�^�(�:_�[��;��Gݜ}[+NX���9�.l�T۴]��]��$�����rl��2>���ʀ(#�}��N9�z	JڴZi$��O;��ֿ�A�=���2�4҂y��#s�/����r��W(�5v�a��'����I��:ǿ7��kî� W����������]e)���с%���[�if�����i�T����<>=	����MG-�?����l\��@�$�(�F��y'���/L�T7F'�$�RچކDz(���JѴz��Wje�AW�L,��&�E"p9��Ͼ0��C8`�o1����Q���L��@�,�j��r��̭�'k��1���f.��i ���Êʞku��R^#X
���;�݄�b_���H@�D�PB9^q��:SKD�k �N_U@�2���	N[�Y�%.�s�K��	(�������@��-����d0{W1��\�*�%��}`Nmvd7����.3���B����;��Ѽ����Ȃ�WeJu܊�'O��N�ߡ��m�U43�&"�^[������W��D5#�2��!���z�u'��5<���5 ���y��\�v�:_l 6e�7RDJ4֊+8ũ�Q����a���hB��0�"�dX�v��N�p�S��p{]Q�\n�ͬ�H�:l�Y=\�F$! ���`��h�#��^$ჼ��NuoQ��ϟM��  |��v�D`�E���;�u�;���ٍ�Fpdʡ"�Zv�\��B<b4ZQC*[�Zp[f|��N��G5��Z�١T+4��M�G$a�� EW���̾����gѪ�Q�ܬ~���;LR��1B�VБ�)L��_����s��*�c��q�+����m��bՏ�z���ۊ�p�a�:���Z9׋:^�#��$E�F=]Tw_v��2/�ʥ���R�xCo19@���%Y�!U�{��A�{Wa�����3�C�3����F7���t��\��j2�r��$�BZt��'g��}�!���#�#ұ8p\�[��B���Ȃ-X�ނ���v�.��a�ǃ����v5%�BY�����-�w���4�e�6	�ij\��]4ǊZR�l���K�w�f9���D-���SKϠ�����H��՟���}����u�9Ж��E�����e���̔9����cx*����_��v^kS�;�RM�d���X���M���:��/
��|K����2܎�/2$a��x]�z��ҋ���-a�!��40��*R:�rGnQ6ꇪ�{`�ڻ��(��<.MEqm�z�gRF����e`�9�̓_�������|������^�h>�5��׻zt�ےvU��'U����C������K��UG*�mїh�����ƈ7H�I�4i�pϗS^ҝ�+�&��N�!�z�k1�H�V��Uv<�z@����*��� ���B����Y�����QZ�7j!�S�+,�^V�e�
~b?Ǳf3G�F#/iz&�Qxb"�&K]�!/8�~���\���a���-A�GW)tb^g;�[��\<�!\1aɧ�.$���������^x�S��$a���ۚ��x��h��ac�4Ƴ�ڙ�0�,�B�[���<
HzS%�� �2��9ۧx������X�m�i5���WA$�����izuw���T���ض&�ń�����������pRI��҅��!^����L�1��5s��ƨv�<�<�1hJӼ�>i�A��i����wzŷ�Y�è�:�4�Z9^�p0}G4�H��� ̧y霤n��5~�MhK-j��|Jz�2Ā�ew�ĳa4�U��������(d��Q�������W� <�L�5����uq%��o|�'|#M|�=q�������i5dW�}#��v7�� _���@���¹#�z��b��>(�a9�+���)�o�����?����X'�`�'(��n����Ԑ�5o��5^��ژ�i�]wJ,��1L���2��L��X;��/3y�u�\z]�f[H�8}bEq�m���<���A1ȯ������v�h&��ں�ʘ :f�D�l��Z� ����|J'�Y�:l�`�$$Ū�ea�j���iA�G�S��G� �\/U4%�R�ϊ���!����=�}� ��C�ʚ��ɿ��\�>�Ӻ� %�:�s5m�)��X����>�? !�lmC�s
nG\�
Wي4�)��o\H��
y�%��?nQ��>�^Z��*��$ ���h�E��_VTpa�W�F24� �=ֈzf` ���G�uu�na_�f�b�9l��H��c�1#G�C?Q�A{i���9�F�2>3�u����X�o9#����{���!0�D�D�a�dWɂ\�Aa��[}�R�IV5Q�(ӗ��,��{)�^��
x@�}�Ew���=�"
z�� T�1:T��U��Y��Fa|�KEiPqw�:�λ��K�)r�M�o�"����mGݕ�K��ȒΊ���vb���\�lVYB4V�#�;�m�+2(.��y
�e�Z7dMn|�ٜe�Lr����p&�mZ���n
��|�אc_\6X�����+vVU#w²����$�ʰ_
���9MBк��DR!�g�v��@�	bk��D`|U��]�k�]��,��. P/q�O*��8��b��̫��;�g�����(Kn'� ��W�֧b
ޝ[��Cj	�D�t����s�4�n_㾬Ů��&Xy3O��s[үK����YW��z��$�	Q����gl{��ZG#��o��e�����a!4�m��u���N&`������ڞ��VQ�����3�X���OgO����!Q��蘥^�)pu)[*%Z�r� �j�+:ݲ������C�g펌tYz�VIɚ��k@����`d�/&EK<�Vi!{�ˢl+!��YU췗q�b��dg>��8�/�أ�6L�>_	�gم�JBV��k��!��}���/CH���͟K��x�iE��U�׫����O~WBT����[���*�A��r�F	�������&N]���>I܇kQQ%G���ZH�T��z����UR�v3�(�	��Y�4���-���y��o�����}��Pø�k��\3�'�/$�C.i���WËz�F��gV؜mg4M5��|UYʞ�=�X��� qvֲ�=pl7{3����/��D��ŰJ]}�8����劏p��N�mLI�|�5�MK-�$7yO!Y��@�xa��V~[Q���w�5 �\hM�ȹI��

Ӯ��C��������Ky�+��(	*�. U�B�kU������9��o�QLn+��r�CS���� uwqd��/�7���m7����
>\���PT*�X��x�HB�
T�9��!84X-H����q����m��G���]� ���?�5��>zЪ�|�%
$#x�4t=��e�O�!�)�F�l~�G?�`� <�@����ڷV��
˸!H�������;.����EoF��{����Y>��j�$d���Z��^���m�;%�z�sp�����-R�+ԁ\㊆�2eX7�OFЏ�����|9��!1˿�-B��&��8p���b�<,�{�1ni&�1ٳ�1�
�q$�:�Ǐ���j���[���vC1翽��Vi�I�^A�CEC�s�As��t�Sǻ��k]!���y��ʫzj9^�� X�/���-Igw
�mF6{��y�ߟ�n���F�������$X�'C��������df�p~�Bg.���M24ۙ���J�f`�XwBƥ℃�!4&�"�f�5�����N��Ke_����ӏ)4��GW���*m��dj��G̻��h����P�)� 4DU4-����ƀrd��oV@���'Mw�䊓8�9>teA�K�X����?SN�� w!9\8B���x2�z	轭N�n԰�/y� ~��h��gn�:�x �Ć�����P1�����[Xv9����{��Q�����,�3��e,U�3Q�������@8�r��ȓ�fW�37��	��n�+Ԗ7�4�f���):Y>5w��`
���kͧu��F.aS�_�������1�᮱=�C!O@4Ws��!���9HY=�x���oJfHH\,�t��;�qM��Z�G~�Upog�Ξ�G*ū���7�:G��e;y��L0!f��T�xr�s2����u7�V�ƑwFCX��}Dap�y�h�c*�t��+���R� �T�sý�,���z\,[x�����Q�����S _����(��-�)_Bbܳ?D�uG�p�:��g�B���4t&7�5�6,�8q���WĞB]Y���_k�J/�ӭ�n����jm���4Q�M���j����W�`r��A$�j9�� ˓3��(�T{J��.l߯�ND���c��O���I������x
���w�Ha�39�Az����,cԤZ���B}�# �#�m���n�x��q�KQ:w����|�)��ŧ�#7�=ɖ'�s������=5�WH_y	�/��Y�a.+<s��h_�b�Y�`�o��u�ZM�I�С���e�c�yV��� ��ϩ�LS�r�V�`�`%�c�nz���渰]�+�/�{)��p�0<Z|��1.���4�>�\���$��WXA=�]��CE:�D�"47�0w�kQeI�f'���Jێ�X��Ţj2��&�n���$:Ɉ���!튫,A8-a�3�t_^�E2W���%�Ӛ9�����\zr��<��2pыv]aV�H��x9G}a8}"��������%��8��a�GV���ץ��w���u��i"�@���?�4'��^�p�a�,C.&c��� ^f�@h~b�)��Q�sǡZye%�?Ğp�0��P�?~� �x�iٺ�)���iS�/�!�j���̤��磏눎�
w�
�D!Y�h�m]uͪ���ɠq�u<�,�\v˽�]t�Ϙ��dc��V]��
st�g�\3OY}���!�V�����y�S�|}����&}��E6���b"���ܻ`R��ouy���K*����Zl�1�LA0{�"AX�%w�K~1���pM�����Tzcr��&��Gڣ���K���	>B疟��h��P����o���;T3��+�1���^��$AB	�<�x:�[�
⧊+�7M�+e�S��P���r�$��R��Lm`hb.��__wF~MVs��-��pw�!�o.��8/��v-�%��ۋ�%�M��V��,2��X�$2��p�^E><�{�)�H�&�2�h�F��Y5��;�J�U��D��UhL���#�X�V�i+#{{=vQ ��U���_Q:��zFW���։]4��̑���F�����gaRY�u/�G�%��n�f�v#N=/�`s�����6���{����
�$���������R%KbuN��T��{y}�L�?����sI�]�zn��Ϧ�4�G>ĉ=Y/�� {[�"|�/��_H�lp�+���Oӵ� ��G���6�+L���+����l�Ht����U�P~	�U-���HWK�E��])S'��[}?�;��bWn5�`FYN*h�Е���ǂ�����L�������xQ
H�c�	�D����t +�]YV��Ԙ�"���o9F!8`5h�;0�I���6��P�UO���g��o�Q3��u�N����ݍS�N����gH}�IBX�An"�v��)Õ����Vm�h�{c�)K���n�1� �6"�or�r{S��i�Q#X���o04�γ<kD�{'C<֦�����9��g����������e(:	!�?A�H*c������p�Kj�o���.�(a[`h[�|�C֜�[��+��(���\����	S��ap����E����V���KT>�=[w6]v������٬Z�oҚ��g;2xr�r��2�,P�z�������q��|iZ�����&�9*�ӊ��t	Dۤ߉!���q���Rg\��l���l&v�n�]��Pn՛%.�U� ����%�j��)n�9a��nL"Oá�3��CE�j���
D�Em����Ri��uT��|�x]�RO="~W���ˌO�A��K6�5�2��.�hiå&��f�Mg���(��; V�d�qy��J;�zn�T-�
壍�ͪ`Ki�D��e*��m�2�_kδ�E �H6�'X2��5�5c=�Q�A��nI�t�����v@=�~ �nvDN\Y�i���9&�!���7?�a5*s_2w�y�Y�-ƭ�D����|����-Ҩ�S�ѷr[���y�l�T'��P�Wq�#� <��M���
���Y'̰�{�+�v��&�>�yLr���E�����q����G-2�=�?r�G9��pTq͑
�ǀ��`��l�R��YL�i%��V���gKs:�O���9,�Rm�|7��Һ�N�9��az��Ƭ��E7��j�����/ҟ�z@z�m!�Z���|�=��A2z;��aFH������n@�������NHn&�c����Ü����e;X�i�l�m���J����2"���|�c���ƿ^�9�F����"T��#�C[sIP������Ŝ�l�lu��
x�L~�g�K=*,̏��f��Y�TܿYM3S����#�Sl��w�:�0E_���5Z��=h:��hn�&8R��%s��x^�a���!��6�d����-dJCKl�A��-Ɯ�([^&[��HJ'�{�"�N���=\@g�O��b(�=NP��HOi���\�U��L� e�6�������R\&_���*��H'	��y�`���axe�'ų�Z�|1��BǬR,[�4�e���+w�TJ� �����U�4>�B�$�t�R�N����@���|�j�kW:.��Ɠʷ�I>i���~�L�y&�����TmrG(�xDe�)��(�%��x�*��@��k)>���}�U�^��eEm��*��-�X�ņ�z@��0���ƚ7췗�9�&��^�iw�Z���XUxK��k}yDW�.�;��9+�3���r�i��E�#�)���SL$p:$1�觕j���l��a0qh��^O^=��X��׋�_^Z�����۳���ZGd�j�#�B0�}��Dp,�_��� ,�s+���,!?�cpen/�Z;U�b�_y�Rŝܻ�������O.�xxF���|�1i.�kc�!%@�Djx7{��Nh�2fm��c��x>)�j��	�&o���\����ȇ�="�+���r���?}q�譚�ܡ�����peX��*�YD�`��m?�5��`��$�	 ���i��<Y�u�1�����^�=�r!�1��8m��֧���`l�Dt[�*��6߯#)��"��hF����+V�T-?�M����AbRO��O�1��Y�X\0�JA���2P�0Am�B�F�Z��
��+��O,�V�X*7�e�iW�*\��$X[�Pm~v����s��	�*���D�3�O���h�գ���}R�^����K�e�pۄ&(/$����H�4<�h:��+Lk�ig CX�2%� �Sf��HW�a�E��Η.sؑ�V����Z�R���;�j5�j7�4�y\w�)ࢴ�z�QT׽&E~}}Ā��y�>�y��M�%}���h���0��vd@�~t�+���[Z8Z6F��jEJ�@eP�pU]�C���+�@~2�T����ɯ��1� ��(��4���5��9�0z=0�Ǻb{����e�>��V�y�kƼ/�a�����D����Gy�����G���^����'Oǂ]�2��?jHg�E�_�^������L�g��;^�	g��s�?�m�v'�?�4�<}R��^��9>���@K��ܸ��-gC���Eܟz;A�Φo�qC\C����G����8be8w(�Uut��n�*�x��#�e�
��{�=!��&���?�HB�4�a!�����h$@`�|%d$4j������ݾcX=���I�k�ߑs�c�D_T� ����b���J�pX����ׂ���XV�u�nR�y�CQ�h�Lr�t7�ےg)�:�.	���k��\yj�o��Zf�:0�1u����TѲ��y�=+������9��ſ�ߠ�.��Ur���6�7�n:���?-����AAQ	"�Q�E�����8Kd����X�?s7δ9����X�Y�Df}$�=+�w��^=��%P��N���>#����@@˥]�*��wϛ����D�q���O#��������E��b�"X�*0��s�.���e7�����b|��s�9	�nG�����2�`y���ХT���������S��{����L�˧p�A��c���só8ܿs��Xto���A�J[3c�<CS�	��X ��ę&�k�~��]�%���
4q�����eoXT�
,�ء��w�S׋���gl8k��Q2�O�5�3���_�J�뗯ԩ����(=`@�#R��]��!�s|�]f�n#�VB���#��D�`�|j"�+�R��������q5�"G|T�Ku�<E��CN�Y �a=<ۈI��2`����9�8�B��TFd����P\'4#�~���U=2������W�D�,Yw�K��Rǫ#���^R�f,����y�C�K���{����-���λ����b��p+�&������F�Y'r,�g!k�^��N���і�����zcL��ӽ�����'����_�Ľ�$��7��n_�CߺE�D0M���Z@r|���g<�4g�N�J�T[4� K���Ĳ�2�W�u�pz!����J	tS�TO�ڙ� �
s����S���~�	kSƂ��������͡~���Ӳ�f
f���{g���\�k����畜ڭ�絼�_��/<X9	7N�	��Y8��W� [:�%1o:��9��.�zp�7�.>�+w�;�:|T�q�C���`�-!W�'	=(�w,�O�1���̴�"�'���h�f�p���W䳌W��5eI� ����e�J��<����ݷ
j_�)���ٟZ��*�d�Z�7Y�+�T���Q��*rD��g<d���X��#Z�w��o96����=9���^ty�s���8c�Na���đ���	�p�.���:^y��MVl��P�w�J�Y�tC�ښҜ�1c]�������U
Ld#TP�ZDg���9���삟�5_�[���O��B���z�U�����k���6_�w��I��r`���#��C� =D�q���V�e�{a|g��9���]5��Â�1���|as)Җ1�f��_�YT\�wM��p�O���G�St�����
HsQϭ�{\�gD�Z�sA�$R�em��~�������`�O�>'�a�j�=���?5Q�9��7�g�`m�}���@ؙwֻ��y-������	���A���Qx
$�K\8�OP�l�����f�R�Ш��0g?Y�k�DZ�3g��.2�Z�W����W�ā����.�_�'��cNɖD��=�M���aZ|�C[�O�Q���Z�᳞)���W2��1s����e,��!��H%��ܟ�t���� c狰��=��U D�|_����q9���9����oqW>����TU;CW��C��uAme��Y���(��K�(Plv+T���@�rպ�\��x6���'�/<��^ �o'P��3FXD �e1��d-���ȔѲ��� �+m���;Y���гj�� m���0�S�i��� �_��f��o���
�'γ�<h	�ʈn�©׮X��pSu!/Wo]"�H��z��[{P�"�`^w�'_�Fq�e�{}8��k�j�Y9����-��Q]I����c�KN��DW5B�����w`�}�Q��60�O#lHD��WI�^�0�-��Hu�RTW�^��p#���<K�v~�@�f�j�׬Օ1�z2'7�fr{18�.�p�ܖ��6������C�v�
���P.�}?o.Ad7�	O%��0�z�t�u��!��(�#��Fo�Zc��H���(��}�-��g��EyTν{���	e|e��+��H@��佬�(?��>���*K���vl��ð�^,8ı�Yg��<d��>YE!�'p�"��M�
��#� �hs�����n��*w0A��.��������:#�!׶
��DNr��o>�}1���q�!��p+y�>�F��&ꤑ]�
�[�W!4XXDt]f�c}�����N1~�9X�f��ElY(�2k��;��{�G�65;�QN<�1��!x��xRɨ������f��5��)0�.O�d�ڊ��~}����$��h��:&n�D�y2�!�P��&���5�#�\WC/�.��}��S�i4U�����`ё|�3P���X�B1�K1|ͽc<���eN3��#���uy�%#�&ź���$EL|>g��:ps�����E�k�5�b���ƶ�9��F��>ku�
�D��� ��l�$�2�wE�����m�֤��{m�.��&�]�ĤM�~�Ƙ�o4����[�+����Q�N[O�߀��w8��[�0��A�˽�Jf!�oӝDT/�ʫ��U �n������4�7��tf�5HYR�I�,�0�K�8�u(]���.�3�'p)3�
b�0��`��C�?�����s߻&�&0��řK�S<U�F�����eA*_��)?�Hr�D'o�J�[	��^��(?���#��$cM7?���s.v�d���<[���S��n��!��]����\ZRj�+u3[���9�Xۍ��Ό訞[��[���B���l�2��ߜ�@�B����qj��ϡ���[��hm>�O��ԑ�q��SD��	��I֧i��ɗ�b"+?�y8W�)K��[��F�~t_�[�Fp�8^�[&�S��i�N2�S��rxX͊�c�C敔�'��YH��S}����k<�y/v����,��}d��T�d��8���L0fwe�`�g��G*��M�ߦd@M���L[�i�s)3�@:��3Qӭ]��Ke68+7 ���mn��#���G�?�3=��;LG�w�Ĉ��z*+I��u0:E�$Gp�!ߎ��%��Zޖ��jkx�0�"w�����=:{���
�� �?�}�dB$y:M�G�WQw��5�W�D�
 � �4Z�چ�c���F¾>?��Sǽ�gz4T��)����&��5Rq�j7F��y��]-�r����i�#�+�vh��읮���'���W"uS���6$�Г�F������Yo���25��P��y���RPm������=Hw���UU<�a��r��S2�8X����;�8ݚh��Z��4��݈5i{>W��jdۻ~�jeCeS�W�����=^-�����uVADJ�>�C�ֳ\t0c��`:��t�� $��$��E���<��k�4������"4�� ��3%��NFB�I�S����[�8�}��}���dW7���re�1���:uV��Tr*�k���
�.NN��M����K�A��1y\��X�4G;�^ k�n���};�����7-93Փ�U2��ڽq.7���kr���N>R�P��ӓ�y����*�!.���;��}�5��h������cb�)���Zz~�!��>%�8������"� |��"v���ǱD�lg3��R�X�C�C��/ji�pS	!JQMhh����)V�
f�R�#��4U�ϖ[���k/��y���3�s*������;ʜ1�e�g3e!�����2������:�	�e�pf��&���z����1�"�]I 1�6϶Ty�PDQao����n*X�oju%����o#WP8����,$qd7��������ڍdj�YA::��&g�L��:������������+����A^FT�t��Z�j�8��u�eE�;�ݐ��4^.�x	.?k�
���6|D���`�c@ӡ���tݩbe2���i_��}��tm76n",�p
��Cj�@ʎ�W�a<�p7�xi��~YO�i�U�'"����ǰ�o��$�;�L$�z�Oawxox$��h9��OÏ4%��{��K��������~Y�f>��G;������2 �w�����8���"��x��z1/�02����/�I��JO�k*�$�L�6hj�=S���OPC��>a�jf���߅5O��X����1��,>n���c���0wc�
_�R����j��7*4Qճ�d�����]�t���O"���,)�i��_��J��irH~��6]:��*u�M�!0<i��M�;����ޟ���,���z�#��N��T��]�Ó�J��=6D��
��D� \+	��Z�yյG ~�ٮ��Wj�	%'_�ϣ������'�|si;E��)}�Q����&^�N�W`D��G�7��Ko�'��O�*��Œ͘b F�x�cT�}�Enp[A�5�=r=�{�z������+?�ɡO$��<�X�dR�h�%�������#�&U'��`}f5��d�V����Ҹ��vy�$o�M��o�t�/�0�'��!m 0��c�쑬4}��K�ؒ�e6��(Z�v4#fE���Mtf�0��TJ|����B�U���#'C��ڪ90�	��������!l� q
)C�O��Z(�?Gn�J�U�"�:��U���Z#������9J<�8a�����`�1]��q3z�u4x����ss1�fbzH����9����f�&�\�����"���.?�O�n��XB�=p��دq)���(�睑8vm4l3 ۾	
��'�Q&��`	mmt�Nj9���̵� ���ݼ*��Z�U�Q�yg[�� �F�A��Y�ǒHF�q�\:8�Ǿ�{^P[V4]	��K�����]�
z�>Z۲)��|�E�� M�L�5M�&#���琊iJ!���W,y��%]Y`q2���C;��,�*���Ь9���y�7bj�2;�W1���]��{��-x�B����U z$����d���I�0^'�yX�b����*��G(�3�O'n��~f{{[�`�21��gc�W�AXc��L⒩�O���\Y�3%O{!�Y��1��)U�㹫�Qu��0)�O�z%�H<{~I3�>���A���y�(��)�@,F�����"j�TD1>*c���Ǭװ?#?U䬵Oq�.�9̃��6D����a�]q���CMD��C�з�}"� �/h�*2����(�X���D%!L�Kca;�<�Y����;@�� ����*UFă�c���i+T�4�C�D�&�١5�q�:�K���2���{�d| b	k�3�u:��Z�92M������C����c�Y�$�1�v��v�^�/$��(���,�M_�1�֜EÚ�f��-�)�b��g�j��S���wh�!7�)����8D�4W�b5:Y� �ӆ�Kf\i��'
�gX6��Í��(�YvT1�wEH���~���1��Pxe_�h��+�z{b뎌I3������ըo�әi���W�&�7m�#u�8���ykC�]z �w�p4�R����=c�GB�L�I�M�����O@'"_��8oRrs`�#�B����nM��0*��[K����F����V,`sX�h/B�
�p�P�S�+'�Ͼ�Dy�\���}k܃����"0�I����ؔr�"QpuPo�����G8�la.c���n"8�6����DOQ[~���M�z�(4��0�1-z��(�WoW���}���\u �����$�2�ryR�����[DQ�%�h��ڿ^U�U�c�rA?�p�H)0��6�,���TQ����6Ak�[��QѴ̮��)nk<�x��1,�3o�j��5�kŦ� ���c\���������1��W�Me9.@zX�<���^vx��-?�h%n#������f�kgnt�;��}����\��rpy�*A��<-�5F�k��H��2����9mΎ���O�R��&s�L+͡=�E�]�VL�ct���PKX*\�����1�@L���1㘾"��D�B�Ȏtb�;�}�Ad�zj�5�գ��m�i�XGܝx�G�����4�p�/xa�Յx��E$���u��7iH����9}��;y-W�P�.�HJ�ǏZ�^ϴ�P��M�d4���D��}&M|��?�*u���,�W/��q*�!uL0��
hi��[]Ku�Bb|�n��VT2�#� �rC��/b��OlP��Q/���I�O��+�9��e?\��y>\J3���X�}�jk�C/�Y��n�nJ#�j��-�"�biNJ��Ա}�P���cx���عʖ�AT(�.���V��R��Фi�a�يH~?i9>8	u��L0�(9ƥv�ݹ��S���<���f`���P.��[h�e}吠�6w�}Kl���?��M��<jr��h�Y�y.￿�Mꬄ*�a7��z���yF�n[Hi5T��L�U�*�_���7�1r�Q��8#X)��n7l�ŕ���w#F�i�P�]nX=���]Ce�kZ�ә�+���ɩ)���BC�@�_	a�#8`��[��K��x�v���v��'$�>�:x��g�7�lm3]e[�L���_���K/��­��v'�8�����5�6��z��u�	��вFAF?�(�"d4,�N>�
�_l3e����C�1����H�,�w~�j)�,s����*ss�s�_�������+I���t��y�t#����K�7�ȅ���Iu��=h�a�rb�UTe�ɉ>�Ұau�ѻVB��j/T�g�uJV,>,�"���.�Fr �$;k�QyQ�e��v�E���0�
���瞙�8�)W���w�gI_�!�z1���
�A�N��o�����W:����e]t{�4	�n.��K��0�N�s���2�¤��촩�Ez�)zwu�������$gAs�>�����*S�?���UĠǙ@�O�qF�o<������/hn�+�s����q[&�ua�\��&���V���BMD'���T��L��u�n/E�e1g��Z\n�wN��Tm�����o9�Ԓ��&H�w�/5��-f\�,�4�1��I#���]��ib�ܧ@��i{���JW@�192D��Y@���g�f6����/8+��m)Ṽ�O=����U׊mR�El��z����|�Hxido��8ډ�#�!E���Ht��lm�?종*�j��]�V-���qL��*��rq�c]|�v�H�P"5�o�y���..z_�ꅙ[�������J��>�N%X#��K�g��>;F�R��S87F8�C��,���]��J�?�+��,�:^-Ƞ��e����$��)��b';aXȏu�MP(=&���$8wU�NTB��S��]����y�瀱N`��w�-X�\��\k�"����]��b��"A�2����r(?_\�5u��֝:���ldO�� ��Wd)1�?�ah[��rTYӀxjy��e�6�rV˞K��Dw�D�d~�/'|.�w����P�������(�K`���!F	)Q���W���d�@��o�8RjŰ�� �qR����yg�	B`ǿ�
��"8,A�#�$�[o�[�tOk}��ry��;� ��`TXP&���!}Q�O{ͦ��5�;�o���Ʃ�K�?�3���p)S�6U}���pP3��K@�E�o�Q)1��~�f٩��dR"�}����>a:o�� ٗ�x�׹�2Y�'��7��j!��{�BE�6"W�B}V�'@�#�e�����>s�C�/タ�$_�f�y^5����kV`�-4�������dd���!K]׾��D7胈����(�� K���8o�L�7�i���v-�2K��Ƕ/�"l�rP��F-"��dBei�ƀl�GH�1����6P$j���o��Vue_�OBl���3��x=��${���'�ߵr�L��mԁ~�}��[����9�Ӊ����&����=�~��s�`H:��c��C�p�d�g�����������aV�����6��uN%'7��ɳ<����e�߸$d�+pp��N��tEܟ`�)��-��y�Qb��kp��Q�Fٍ�Cbhd�|�� ُ8Y�#��c4���2�� _ln�DUI��k��u�%�D�T�g],����P�a/2�/PeAZ�vq:Q8G���k��^0�f�?*��mM�vn�4+PÛ
֥�A�Jt�c"�G�5�j��@�-�2zq2
s3��������鍲��(ޯ�<����aܧ�͢vA�n ����?x��x�z��pp	�._�SC����:Ǘ�^y����-1^�2!&�1���z�p=��1p8h$ ��R^Ti��G�e3��/��O8�)�B,l�Re=�l2Q���d���u���e\[G>n=�g�36�W*P3d�o���p����k��u5~w���s	�Ls{��k�9νw��!'�)��RҴ�*�8k����D�	���������@�y�h�D�Nވd�^Hx���B�v��^�F�S&h��ɩ�C��)ɝxWD�������L��o�&�]���m�t������i��A`�s&�LH��k�Ѯ���7���.��wC������HH��|&�F�!h������_�����|D�%R[������T�y��y.`T^�6��$�Vo7���,�o?�(�n�KA74�i�����=i��'��7����W}��^>&��z(����V�륺��[[<��GCzEx�찳,V���W�a�<�t����0Y�& ���+�L�K��c4ԯB��T�OL��/~G�Ç@է���u�I]}�<��%�cx)(�9�r�.67�Ѻ�na�[�!��m����~� �J0��g�dI��?�x���^���C\�S=<r=E�$�}�菔��F�{쨃��C�4�&,O�4�o�en���E�4��ƁhO�Q��X�� gh2�W�3/`WL�����P������K�8�V�޶M��2��o��ު�t{p^<�~$��o��X�0�L��������65��X�����T��Aj�Q�E��e���;h:T��4!�Q�
kz}r�����AaZwZl�E��b�+�q�stΟF�xJ�+{���i\N��Yk�!��L����]M�g�o�ҭ[��s�&U惠-2�����PRS���b#��)�13){�P�ܭ��C�^��75BB�Ǥ���t� ���*)��Y��A��?Z�%�g������t:Ct)_ ���ژ�P��wH@����87.ۃ4 �@��ɲ���.����J�7�6�ƿd�|3�1��#dn���w�p��ʆ��pΘ�n;��\3.�&��;w)��L�/�\JsҠs�*�P'�5���M)ؗR(:JCas2��&��]����ٯ��o��d��RH6�r�Ĝ:�Xc���'wX��R�:��TBn%��*��7O��-G&��84&*��Ҡ�L�:,d�i�������-)�a��B�}�����۠�I��h����R���)����1F^�e��xp�����[5RE�W���U�&N��'V�h���,�G���MmT��3�gfۮ �wK�.���C[�}�]W��^��GLHd��}Ľ���qw�ߒA�y��<��@���W�|x'�4u��ڱ��T�Ax����!��¨�JR�ᖦ��_���v�ψϹ[�&E��Y�4����ZeP���kb_�=ݲE%P�G�[��˭��>�x�?ww_��^\q鼅˃e,��"P:�>��c����K��&��lf�(J ��TyWv� ��D� 4*$H	�G����?�Ւ�r�����ٖ�oz�`��k�st�8q].���,_��m�<�;���^HfF���"�S�\�0�2����|�C��ז"�i'X��1(�=�Ǯ�|�ld��AHgp�!��AO�o�*7�!+��*F�s��O�7i�>���A���ɸ�F
�(���0|��]pHc���dy�2��߫�~5È��a��H�'W�?S&�2����q:��g@ʜAr��,`1x��������̬�.E};�c���۝YE�> u����pb$� )��}�Kj;�,L<�,<Z�R�DT<^�=�J�*�L����]b[se��l��^�q�����w�q��k�od��W8�F�����n��^$���gW���kT3&��D��;!|� 4+P�Xb��W�g�:e�%�,��8Ct��&���.ٹP7�.�=�0�@o�F��X�^6����CW���H�3BZNA�ý�Ӄ��4�-b#������Qz��Vx���ok +f��ݴ��k�X�dK����n���`о ��U����.�NYZ����S}�k?~j�wKG�����[�KQ[V��������0eZ*^���	UM�:���ש��3{��d=`$s7)~�t^㿪��
����<�(H��: X�"��5�;b)�ÑB�	�M=ED*�j9͊RJ��=�3��B�ֺE]��l8gHwԖ���Ja���xI�cc̶��F\O{ԿA�BѺ�V-��2xߏ�д���I��'a]r��8�|�������"3c\Z
�.���*A��أO�x�p��Mg��vdl.�>:{P�4�R:}Pn[�EK�x����yFp�'�	�X�i�..&�d[u�+\w��jÇyyX�_�7O�k��aRO��>�E�J$ɶE� �f���5�u��T� 	T�9&|��]`q�]�@���������P�@��Lt7�@w�MY���x�e����+3�D\j�����)�#B��ھɒv_̾�1n�C3E�ϕ��Un$r���F�8���dI���b�j^�&��{���@���448z�O>�;:�x�=��
����]�s݀� ��Ή��^��*a.�H��Xm��@�jJ�����d��=�+�>�k�.b�9i���������Vnm�/��?{�3<ŋ(qFϕ�*����� U�\~����[��w{e����OA���ǋ�XJ��!?c��k��V�Z�QC�������R�����b���&��l"xםpwp�rR�����ͭ����&�g͏�l{��`�ԋ~�h�����hY��&�2zL"F@��iW��^��ָ����k�L~^1�6�����Ż��S���/��Cqx��%���/q�!�脟�\�* y��M��ʻIJ~��n��.�a�:�'����!m��^k��s��"�=����i�������%���Ĵ"���وяuRfO�C}��ċ����9<b| �y"Q�Ô3��,f_���o��p%�� >$o��� 5��e��l/���g�x��D���*$���
���j��s�����F<u���}�zX�
w�R*�~�d�WRq�	U��6N�"�Lq�)u~fz�%��5!f�̖�|���"����uo<MM����dK(�'A{g���Wċp�yГn�ȳ�c(��]n�t�[a�
���E�[��m��8��ǂ5�������ڂEM}5ڸ�9"�=�A��¹�S��+e�"�(} �_��i����ô��� �Wo�cp��Fu��?+R�BV0-i�`��8ZN�6�1��e�����ψ>O8�'a�%�w���q|r��������\?^��i��}������'�����1�@����<�Y�<1�N�g;�GS��ʦ�n���������;�i�VdW����x�T�A�����t,�Ȏ����[�v�٢0����'A,��Kd�C7��[�l�����'"��qH���8Vꁺׁ��{��z�ЩG$��{(�kV�b�JA�S8~�q�8!��j�y��KO��s�u05�$��Y����
�v�8���%�v�==I���rFB�N����#�3�.U��6��H�&������mG��Z�y*���URYV7����YA!��u?S(g/j\�pGh/����B�i�!T��'��F���\�x��>�X����h�b3�5���/? M�ϟG	>�ܕ5T�{Öd�x�-�����}y�0j[��x
t�f�qf�d�%Q�[�e��5�ou�"����������C�M��4�_9�r����^c�u��@m���'�����{���k9R'+ʛ:-�� W����[,`4Y�o��B�ז���r��@Rt{Jr"��5��)�zoZ���<�sB��r�Ea��c���$���2�F�l�R����k}1����z�H�h&����N�{^/~�W����M�*�l��d������
ÅT��M�8P	|� �݇����
I��W��R=k��dh�m-�<�w8�N����/\1��#_� ����R~ߕ�E
����E�u}>��l���xml.M��2�ul-ұ.5��ly4D#�R��&m��G�Ӌk�[�~���.�����
��JĂ|�k.��V?s��9���L�`,f��:F�3�x����b��y��Q	��i<���
�T���M���2�N�#�H�շlM����L'�8m^6�ܲ�9��؞��!W����Rȕ,�9C�������i�˪���+?=�7��20m�(�����!ZE�<�qH9(b��g/�7D���*�#�YH�!J��Q�����k�`_'�!���J�-���\��<�3�y�R�+����ES��g�����7c*}�H�~���u�����%�(H�59����T�L������IW��,B�+�lN��dl/�61]�p"[/d2�\�*�2�����{<��iD�@�l|DV<r��L�o.�r?������W��,�'��^���<M��*��]��n�06}I��8�TTR����R\������xC�(��ǭ!��S17Ī�1�D-�C�io2�s�v�c��ėkA�~�]���?A���ɇ�KϕnMu+H�(Xs
�q��1�e@>\�_~��DZ����ro&m ]d���ty���f���=��WS�����`0�/�r�1�5�k�T4��uKNG���=*����O��]IJ�Dšm���|4�R�zD���#`ٓL5�n��_�o.!?��_�`����Ҙ	�&B���N�zd�axm�teR���p��QH:�2�w����oϒ��R�1�X�P	��F#m���BQ��˼?��&��dP+�2�ʯҙ�"��qSSDiUa��[��_o��7H[�@�+�[��{<֜f���F����F�E��M�Nt�Y8��H��P�1x�<.)Ci]�?��Jw����t|#z�h�TS��̙�(�;�Ѯ���^[��q�%Z66�Y���FMKM��o7f�qT���hȰ���$�Ƚ ��5�hm�b�F\�B+��5���fAyJI�-v�T^�-'W[��]+�Y������;>!%��%\�س"V{����3����!����9��y�G<�Q��.����&�)d��~8�cYH�L��?V-���n"�q�^�|��ŅCN�2��"7�Q��6x�R�/R6b���P5��'k�w|�G�7�CBYO�W"f�{������c���~��:7f���@���+�į(Q߷c��'2��D~��&����Oua�I1��w�EǞ�^��ͭ=��wCg�Y,��P���.w��j��Uέ�z��� J�"����zk\4��_�S�{h�NX�iu��M2���^�QGV�-�OSq�bK��Y{Rc0ku�c��k��n8��r���1�	��l��q\�~����2�zC��0xTN��v��,��u��+=lp8�z_�gx&��O������)z�ZT1]1Sr2����� O���k֟͜�괓\�X'Sx��f��57��DR�*�����1����	��D\F�0[X�f�/T�m�ѱ����5{��Z�ւ���a�\���K�ב�������#�����B��;��V
;#/~Сa��R�V�����Gi!�}vC\ϧ�kOT~�:H�&���\rGr"�%kK�����a�9iO��\3K=��Ҥ .
|� 8�r�]�N^����0�a7���U�0�rM^�(7KU��r��%�526D�Y>�1���j��W�����j�t8c��3���(�ϖz)� �T �8���UW��1p����.7(�s_ʉ�rs������>��$�*�KjX�\�ߠ;�;���v�W���e��l,�Jb1�0)~޺�YE�GFP�VU�=��b?߇�U�
}�r�{�S��"^^��t�Gx�t��$C��Թ�ۑA���T�V�U�Uڬ�kfQ�6Ia�1-x)�I]>T#��������rg����{ݑ�X���#�2ɐ�Z��B(Q�eX��}�#wl�I7A#��I�x�r[8� _��s��@��=j�3U�*��6]��v«��7	�s^qC X�:�<:���|��7�z,��oFX��9�z�^���Re#��X�<{��]ٯ=A-��,m�d�����-f�����X9���tKg#�)6�I��;"��=����N���ǰ<���7��c|���Z3P�3UE�����]6P�o���nfbk�������`C�@���	�Ja�I;���yHb��:�Ο�8��ax�$kQ������n9a&��}%�1�㕎H��w�)`V��j�>��VD��S��|�ޥ�d�I��e�>=T��:$�1
6�y���S�3�j���Q��f;a������m�Y���GT���!�^m�OS�p��Dgut�gLf;�����+!OC�0�����^�X��p�=I�T0����n���|9P��#̓�G>��G:򱨐B�a+�&�)�WEZ^/��˚�����EV&.���h"���t j�^%�NӰAh^�tŨ�-��c��0�)�ʨuA_3����0�5R�d�?���rNp��{Pw���r����� (!A<	&�g�iv|1���+��U������TB/�K?��mc���CKXQ	@�,���v���u=�~$*���r2���C��7g��xiժ��`��~��?=X´�~�$�~�Y�@W��m�6�Û9��.���^D��Ci��/·S���ۭ�A�����F���}nV�v\�j��Ҋ��7&��<D�}A��͏qt�@��>�����
u<-�b��7��@2*����h;?I�GN� {��njB{�ky�R�i�V��b�?��߸`�D*��ZZU��ɜ�LȦ��5�a�����g4�.�)O(������x�D5gd�¼���椄��G��qMZ��x�͗M�Y(�����<����?��5�pR��K�j�Z0�H����e|����5�M
�?��J�U�0���貹��Ւ(}�|��V�� ���������**��A׫��X�sZ����^YP�J$y��\��O^��;Yl��zY����{ޓ�`V���N���67���k0�$�T�3�P��ڗ���8 ��� �������5�-|!^"=�-��ݪ��$R�!5ϧ؁g�|y:6�MZT4�_�ʦ_8�Dis)H��j+����`V|����Ibg�[5h����ݭd��H"�t=��-y2��0�Ux��pTWH-��)w/�_����I_�1�n;�'	�1�ˈ���P����_��շ��5��Өp��^pGa,��k�6UoǬMj�5�ȟ���.�x������y���Ҏ@�a�xe���X��	��]n���`@\÷qf,�M��s�dg����X/N<	ۚ��(�S'�t�B̬�
��=�U��0���u�Q�����������¿�u*qЮ���v��o�!��943i1r�F��5�����H��6��1���?3�GW��[�#� o4�J�����8Ｓ�!�����&�MBe+�~�/
Gd�r"��7�W���!�[u��;c�̨CG�ߎ��=�ZB�實����K;����@�ԯg-J����xe����!������SP|:����
�������O�p0��վ)T�f��`��T�q�����z�mPv���j�(!if�-Ls�8�G��n��8U�	 �3=�E�g �Ϻ��&� �>�]c��`�b_�h����I����fi[,r,5�yݜ�;[O�?��
��Mz_�O�AF��P7/�����>��t҂u��VN%8�?�TG�>��mAg�jw�9�#�>���77m�Ì-ɧ}��&�n̎��z���+�g�V	w���d�-�,"/���J׹���I�#�8��PP��w�Q�{�0Y"T�����uOISE�
�� �28�;E���'���8���Y��Q�,)���'�zwiG��nദ��+Er{�5a#��;��1�b��ܚ�\�/�a� �ER�+ӑX����^�#�P��I�]>s+��v��]?��l^�7m���Y"���39�Ir{��L�\m�W��\��"�6�����7%/�@�@>n��T��6 ��>�0�}ێ�	����hgR�L��f��ZF��U�)"0���̚�a�� ���4�;* �L:-ض�f���_��e�`i$+YŎ���-1" -U�X�:9�D�A�h!6Y`�E�]x6 �W{}H�WZ<;9k�� ���Ȩ��a͗&)B'�'D����ޙeJ�Jh��-�V�%2�v�;�Z5�WԾ��Y��a�8�ӯ���lF�q��2�CQ�,��J��i-y�&o�]'��M �&?��_z�֤;"=�giؗ􄸞��?2�@J�V������k�^���^k%K��K���q���{>A�����+�:V�����_�~�g%:�sL�����b��K�����A�)oH����_��C���R�h�����4q�"�㩺���P|��=_���0|�S"z8�Ŕ�uI��sS����Ѱ�av�[}���s�V^�*�5�0����w҈�h'7��|a���"܈���?et���kG:�5��}6��<N����r��:V�K���Y�w��B�2:���  �2ǲ�6��G���{�'@�s'�r�[���3lo1�ߪ�Q^G�,�r	�Em8y��)�G"��2� 9���P�W�i�{���{Kg4�p�J6�JS�4"�M��]��_����V���J�V8|�v�@�8z��������=t},�@�^�,^0��=g��*����N�:�N�bg�x
�B*zK�N��Gy�&�"j@]ݿx�u����oH���w��~~$ .��ڋ��̤dǩH��{��5n`�zfY�)�^g	�����n�M�����x[0Ayˍߟ���%�g�6��*]Q�20�w�U�?��v�c�?S�O�U
�M3Iz}�g����*�|z"��S��ɎF����Hl�1-�G�O�Eǋ�DCiD��w;��[��ɶ����O�g�jI<l'���//�}::>r����B-!���Z�a9��!5�Ja	N#:������D�6ԡ��K���.<kS&?2^+�|�IH���'������p�X�w��I�,)h�uw��q��t!���7�)Uɛ2;�Y3�a�j�bj{����V�����*���g*�� *&�1��ɿv	��G��}	�b(�'��=+�,��^l��7݄�6e�m���
	k�+���/  j^`�=y_ݨ����>A*��0)��/V��8g�׮Z*�Mz	�m�H%�LŲ�-Ŷ�H�9��|$d>nS����P<�D:�ϸ;s ���wT+�B��>�n���^sP�l�����gFw�B� X#�Ԟ�FՉ�yu�v��JL0�
�,���S�n�t��.ܒ��D����,��S3'���қp��W
�!��yez����vo	%��I���H�g?oJmN$�Ў��0��w�j���ܙ�����qL]��b$�B��G��Q�t2�ڮ�[�_�v�����R`|g�R��B>�l��Q[TJ�*	�4�4q���������[�A��Ր���z�=M��z��S�A)�aďMI�Gq����y����z�����]�G� |8�]Ę�[z
�1��GaS��N:I�u&�#lUQ��? ����KQLO���*�5|�GK~�����"�Ѝb�@A����7�f�c�{�{b�U��]�iߗ���-p(5wW�ݐ>W���b�#7/#du_¾�X�3��g����-�.g"Y�{[�����Rv>���2k��e^���5j��#�z�����oYŘg,?�8���9��s*6w�����pn���9������D�7?��B�C�=�ï&� +�-h���?+�@��K!Q,qЊ豫5�{�#X2���q�.�Ӗ�62ͼSN�a�xl�������U?���7#��)>7�t�R������d�F�Vʗ
$]���1�PN�Mu�J�W���������)`�{w��&>�\z�PU*��]:�$��g��Cc��O�o�H��]C�������ZD�t�f����x&X\�������=ԡ��Wq!���sՑ����[ΘZ�܃l����^�|�I,�I(�o��������E��/��-�Le�=�y����b�@�$�A{2 əZ[��R�;�9�9����Ǻ�mS~|k+R�N̮�ʹ���lq5��*���;+�#���P\������y{���N�ږd�dל���S��$АՖ�{��ʂ��.�A�Bi�Sn���O�%��u���.�6��I�H�?�h�u�I��dFwl�]~}T�`�!W�"v�j�[��]��H!`]�y�� �ෞ�%^����;ךwY���H�����������(�VMQ�BkB�|�%`m���E>��l9z;	*+�,��n� ��G�h�-�� �`�3���=��kYV(�#�E𕯭�`t�v��Q�\d;�m�[�y����2/�|)�ɻ�����"�SZSr �݀eWv�@jM�Q#s�;�_.��eFQ=�����;�إ�r��,Y%}�iSf�p��=��0�F��ӊ��o���?
��`B:�'Ȑ�Bc�����#�[��ú٦��܎���^!I�i?�m�"��*�>C�v��-C�����&�t�)*t�J��9�j�c�Cy:21���SϤ��걲�3C]qk&-������U(m�l$Xݪp�2PVUW��f��* li����&~?B����"�ı���?$�Ɇ���95;��7�۬z��7�m,� ������(H�|�=�9�ť;
u]����Q�#��g�r���ڢ�c�ׁ�+�Ƽ$��1/t�a��\\�:�z6/�a� �4_�������^v�|�굴%P_�?s �V1��X-S�-����2z:Tyg�jf%�H�����5�q
7�-c�NMm����+ ���N��=/%V~4�s�����3�#��_d�z�8B���6�r�:2�ԅ��v!��N6:,{��jP�_�h�l������?)&�TܭIٞS9~0`@O�C��H����Ԗ}�64�6.�L���_z����'�r0t��9P*d��������
&�X�����:~@����g��,�L�fGN�gJ��!����_��j�R�(��q�JjH�s��^�60x��A���N�i�s��1gTV��,����/
��p��w�T
�ɟ{���a*#����\ш���IP��'5�O��;Dؖh&���5��+C,�)����>lгN�>jZPZJg�⋃����J�k��{Cx�J�`5+^���k�"�#[�h� <;�g!�i��o��AC�P!N�b�Nf�,��������"��:�����E(���.��v ��Q��a#R�
31���T��<:��C��MJ�b�H�DY��"�n�k����y��������2Jb/��؝}�鶟��6
��Cz!Ŭ���g���i#X:#k�i╻��})(�b(2A�h����R.^ڀP�P/�l�{��6��$�7(�E��f�3��T�������5t0��8\����W@l��/�L��1���Q���yF���Z��}�^��x��"Z�h \������qk�b���S{���b=iSe����.P�g�Z���(��@|��|��T<�3Z/�b~_��=�Α�}���\�o�?�u�NH��8������mPo|�����v�}�@��� �T��������j�Ht��b�:�����
�[LB����ba��e�̓�0~���2�v����4/b٬n�:�_@���;B��ʢ��@J��^�T=p�l�W����Ll{��1�E���H�d�y�������f<�i�G�
8�@���)�Z�y�O�>`�)6�@Y�-����,'����A�3�x��B��Ȳ�{gt=oX��Jvp������fx�k�{վTCJc�W�!>�w�{�� +_6�#���
Q�>�kL�����K�Oz�����D��BӅP�xTi{�Y"e������Ӕ��-�|�!�8카�Z܀e��r�c�}lEbx�iOS�c�y��h�[�0��4O~Y��K�p�Gl�카��E�A���90&�5��|�2���J�t���KEOwS��J������@�TR�K8���P�`�=�����i�&��}1��w���K��/�)���6ktύO].`>�!�2�&EQ��d8�lq��?�A�\�d���p����r
���`�4`��������x`:ϔo2��`��Xe�sM�ȵƛ���qqw*�T�ƗFxg�Y�����,�r���b-��n��Ř���SN]��B��A�O��*i$�u:J+�?�EHi��f�f���mK��F�O��En8l���D�b���. �s���{@�=I�h�t�x�]^Q��<�����4�M�hS��ǟ˪��P�]A��B?�}���	ryک=��4���~'e2B�?���SpĚ�*ee�\D�����L=�J6z�����[�+�d��mU-� �
�';�EO�:W��F�R^)��,�r�v}=��ƛ/������e��T,;#3Vr��4�dt��.����e��f�:z��4w%�`����Hfy�$�t��<`r*s�P�2W�m^�Aߕ���z����i^�|�WUƻ7,�T���O���.�u@b5��^�XTe3�U��Z�jG/��W�vׁ����o�>�(��8�sn6�B:�`i<�GDH�L�uy��=?�
 oj�&g�pVخ��B-���z|r��U�y��{�Mm���
�Ekn5�;B����9CЛ
�`����r;/r˝˱�[��A���p��
b��Y�/�ƨ�}���D�+����~�Hh�#���XpR$P�P��9�a
��t����0��Nmi���_p2376�i�d�,[KO�ڪ�D�~νp�aj�
���(�7�A率��[ F}���[�lo8����I�AԖ����
Ds|_�)|j�!�+����Y��	�3M�ItXX�G�Fx�#~#Nq"���� �<�lh����W &}8��F��5��L���(�8?��^�m���02����a0rb1Қl���F8�\"�Z��Qdg.��Q]���r�H|{�h(AX�a��ƥ#��]��a^.�X�E&\⹡���y��[<�"���vn���Y�o`��1U�ݢ�JSL��U�{�n�Z��M@k�7���`�	��H�k�/����M����������?�zE�Bo�ㄚM@��Hw���w`S݄D�c�+�kK�P�+чh>x���w�q��ɂh�PG.�P(��Jq�&ZBeR����$���X1d*i���.�M �欨Up�<�T�/�Q�3�T
�F�\A|��j_���*pz���}�S`�pt�g����Yg�1�Y��1����_o�_ߟ�C���{;�N{��j�������I#�'JOqr�y%�X�'� �'ƃ�:��@�2:��s`ݫy�o�z�:2$m���y&���"0T���[M�i��@�n�����W����Fg���Vخ�	�^I��^q&u��ξK��u�ђ*��� s�&1�@8�|��[0��*�HX+a��ݎ,Hg<�#Ib�w�%��yUz�2�ET��?A��f������E��>E-��b>��o@�9ު�"�m��(7$�8�t_��=%`��GȓZ���>��Z�����PL A�0N':���1�d�mE�7�C4�u�}��ԫ~@��	��J��a�w׫�.8١������'���)aM���l�qh��I�cML#l��ǽv)���>�T
hW!-Jխ���M�4��7fxRHOoKR��t.�����e|����J���D'�Ƀ�C#X*}�U����ҧ��4��q�i%��BjY�q_���b���^|�s|���M�B�w�I��$T�l9����Fd��&������C��+e���7)m�6H���|�,��5g:�-�F�|JO���!�d��G&�G��O
_�1C�j�?#�יC0���yllІ���ҕ�����LE
���p9T�D�����ErN�_�� Ui*�z!%bC����
�q�_f��"��&�Sr@�<.�<|G:!�*�D��a%j�aPӦ3+��So�i�.gɒmպl��F,�C�Pap�A[��'4Ѐ�1�u��\�ؙ�(��ZjGՎT��A�$	����kKc^%:��R�H���t+�in���N����,4���i�9�'yt�%҃�+xy�2_��̝\��צK7K���⣁��O�����al�G/wz�+�7��s=�ͨMt�*��]�J��k{--T�[������Dϋǭ��lh�G!`4Fq�
?�D� ��rڽ �&��f<�[�t�V�|vu�ݽ��@���a�L��9tq1�`��"�q����*:��7Hue�S/��m2��@��7�e������@tO"Q QL�Y���:��O�i���6��0m0�gQ�����S�P�v�0M(6Ź��w���h$Ƨ��Ihl;�e���"J������{Cx�'��C�X��	DЇE��'x�Oy���J��P�����XP�]��*h
�s$�W��N?~�J���Ff�ο ��i�Բ�>�E�|(bRP}�/����]����	��k���;-���"֚�}fS<��M���9�h��[�bdk�`�� I$���̵ݓ^UW��=MA锜�S�J���tX*��37Ci��&�s}���FVJn�eqb�}x��h���S���oO!�J�V[ϒ��F��l�@y�P���vJ<��c{��^&�֥h��.�:�����cۇ;�h4�i|lؑ"��h���7�da���4�t�/K��pq"�D����'��������糿�M���hzW�
�opΊ��X��=�/}������m�bF*�GH�r�]�.��Ew?��4� nоgWl�	.X�$�t[�v��"fc�f��eJ_��?�<���C�K �޿��Núr�tN���X�;w�f�8e��I����C*��e����WF�e�p떦�N
�G��)L<| ?P\�lI�_�	�f��}���k�u=��t�&[��ͭ9_��m)9�m���-h���xJ�����tj�%�U���ō�.:���ϡ����ݢD���g!�Y��Ű�N�n'�e�S�
L�d�����*�����g�nai����A�eQ#����8�d �*	�f�kEɇ�����fjԖty��g��з41�-��o����Z;ƣ��M���5Y%�t9 �����%�0� �������|t8V�hBΧm�����`���J_�uS2�Q�nϴ49�c�����Ap�����"�x��u�Ы6�B���(��O�W��!��/��3ķA����C튄ʃ!����W�L}A��텐�oX���=q\G��b=M��A�a���ɺqVV�G8�@3P\~� ��i��c�rS8�m�֝5���g��צh�?��������Z��4F:3���:kt�*��e�s*W��9L��U��"rA�<V�W6��?*2&�σ8��(v
�,�f����s8��ͣ������I��_əYid���A|��W6�'���7l���:���X�Xs�`��KD�㸬�����,�=��]s����y!۬O�,;t��9���j/�jP����]ǥ���0�Yj����Y�c�w��� ��۩j��p��c�~�ƈz��'*� �&�(�'��2\�,່͆�wqe�3��ۃ�������w��� d� <t�ᵉ�)���d��R�k��*���8W�H�ʓXѸ����8v.��cp�;PI�FD�����̲]�	�LA��Zsp�y���o��h��	 ����y�0�?7s�g��ڝ�%���Z�1Z\�[�/[B�0�����+�.� _Ur�Y@�U�7^J���R��mD�E�Bcƽ1_CR��lu��-�"|��m��Vo:j��&w*2z��w��Mcw"@CL\g��D�Ѷ�q&!f�O�u�G���48;k���L��V�U/�I�C�afQ��)(P_uh�ndH�����""uT������aĦ?��n/4=o�˻1ί� �!2�9�n}�����������dR��e�EK"=P�K�4*�Q�W$ɪ�6��v��$Ѣ�^y5��5�0�YG�4J�j_;E4e`��Z�e�g ���i��{���1�f9Ra��ƐG�$.c�Ruv4ר>��%��� 7xF�]��׫*\[��=�g72��
�'쎻��ߴ�. �6�PE�^��6 |#/-����Z���l��Q��a����x]�;���M�J�z�{��n�O�v�]	.oP�L��������� ��g��2�g�_�.�(J�(D��;�w�qZ���H/?X�c׺��Hh���_o�a�,�_�<,9�c�	aF������332����>+i-[Va��M���iӈC���h%T�`/��eCrT *�*�MTo��U{�D�bCX!��Z:�A�Yy����QX���>b�p��Qhk9$���%��'��W�u���A�,�guϵ�D���Q�����kϡ����/A4�u~Fbqcч�|�æ��U6�Eb�Q+G���E��e��sO�I���J�K�|�ȼ�ܗ�� �R���Di��b��y9k�28K"3���.���n�C�O<0�/#����Z*��
[�k�Ў0:z�/[��@�in :����o�ڸ��G=����?w6w��X�F�,�S�i�%�%���/UF�E��|^��+����h, ����X���h�ڑ�W�Z�=�߾�����c%o����:���АBu�Ob>e���utދ��$<��o���X�"���A[�d������ᮖV��İ<�q[��D]o>����a�+���WI�"T�e>�1_��p�[0�m��7�l�����쟐gݺ�į����	?�%�Ý��ݾ�VK���k^E�����HgG��@�n/r�90Q���*�D��/�(͢흀��W��;�b�����ǻ�a��+G.�_���>
���1�Ju��/-��ȥ������8��~��$��"�< ܜQG���H!��0��-�	�,���#�1��с�0
1�*�*��;o�E��6��A��ך.�5��y�X�`����*��F�����x2�׷t�iQܣ�Zܪ[0����}|8���T,��,�vp�Mẕm����� 1�;�ͣ�$ɺ�v�[eMN��~/��
�������$�u�I]ꘉ�¶AH�޺ȡ�3m�B�+����=hV�A����W砿f��Rq�|3ͱK�O{Oֵ��+B�?6�Bt��J���G�4���@��!�rٻ�2�~#�:�P2<K��,���)��}��� i�A��@#�x�<u~�N�^��
������Տ�b;�䓐�j�w��o�ƈd�ЪcҮ�kK[��{��!�4������'������<}�l��~5.�&T����'j/���B���K�;��o�6���Q.(��o�`Z���Y}���B��kʿ��[ &�ʃE	����Ϋ����Gx���5!>��"(�r����*��4b��߂���\�&*�L<u�)�*}�9������UQR}zR��w�Zb��̣%�ssN|	 %f��ǁ�Ҙ���x�[ɉ���ffŐ�R-��2�?Ly&_��&{��e��<�#�}��� S7��/B⫟0H����ש.oK6znI"p�rm��ђH���XBJlUo6�	��C�8$_[��^���;�bt�/qq)8E�ӎk�~=O}b���� %EP�o�3R�q$��|0��-?n������"�J�9|�1�e>_pe8G��}�E]׊x?����έN h���)��B �X&?7cLn��~JQ�Mjs��+��l���(���ۖ��Ժ��J3�~&8��8(��b�k��r��Q�D.�O�xx��pt�)��G��,�W-��}� ��O��Г�0k�HE7�����y7_\��:��=GC^�����_W�Һ��ʥ�mHI-a@K��'�Va>p��ܣ۟�h����0�2�Aܺ�`
@|��h�����ٽao�ou�nV[~��W����y��R�����my���α�H9NFP{� �� ����)�b{澡T�+���(��\X�'�]�� ���+�\A,_T9��㸈��z��5#~]�d���؀����_��L��X�b�`aM�� ��vհ�������K<�}\0�����!-��a�D�ۄ���R����u��'��,c�W/w�`�z���`8S�[�(��0+֐ϵ�y���WuT�a9F��&;`65��~� ��M��T��W>�*9un�w��
�C:���f��\Oļ�$S�8(�b�2~���[�8ym��!�:L�(�b�����&t�5Vܛo��S:�]�o������n��_��W{�~� iN��>�5F�V���'��d���Zh�2��h�\i���ޖ¿��
��1���KQ%���-Mo���Ec�a2�8�H���3��m��	��WA��'��`�}g�h�D����C��`�.WA��ukr�%���K#̭uX\L5?����~��!�U�/�T����{��~ R���򧓍o=9����ym܈l���\�[?ט����x}��8�CN���#zߞ�.%X;�ad���F��@>X����Һg>u/s���B���<������}V��=q[,�5����w]��'m0�h��c�I�6M�����-�)g:�W��&D^��[V�����V(;qxroL:��/�TN��:�+�S�h���g�l��H�޻+�ȥ�/I�}���`b�+�Ņ��ٕ$��G=9��j��u����vPh_��ou`m;��7I��sg�¦n�)�C8���z�>R�%S�{���C"�nt�ş�]A�~J�+GXR��>�~�
�l��V��(�^���!��8�����������h�B�Z?�������1
/�I`h�&�d/�_��1?\.�Sz���(
�T�#|j�fv"��Uΐ�숁5�3�K��gfgd��Xr5Q��*ss�}���?�_?s��P�{�T]/�K]5��'��5U����oHa��.�����g��)cN��#��� ��b����ַՑ5y����Ss�4 R�Z�}�b5�xa��~;M��{A*�����t�E��o���9��t��s�����Z��
�:�lA���kS^q�g�ߘK���c�4&�]�w���9�^)�5#1�ԙt�]\��|k>:���s���Q��MC�~R�E�A���bH鮌�*b�(���ze��8<��REKG��cj���t4�3���"$֬9x��d����쐘o �r%)�D�<���+�>0!��(N���OD�mz�/E�n_E��ï��oP�F㌲�q�ƍ�����!	\����;?��Koխ�Sg��oP��p��U�y?0�Z�֭$�7P�j%+�����ʇ�e�n]54��R�����c[�}��Ak��������K?�i��̠��~��Zq�̅��a�7����|G���S�}��I��N��29t<�hg�%�@|j`�U�ӂ��鳃#�������.π��}́�\#<�0	�J��c�2�l�޴�����xǫG�+q���X�0ثf��$�����%id�=a�N�4@����S� O��lNӑ�����T�g��[��
%�@�����	�B(�J��~�I�H�͵@	
U	\�|;I~�27u�U� �pv�
�E@�$g��1���թW��u
X�Of�����#��%���9��
](h_G�<D<��/F�,E��X�^��E;�tGHR�	T���u��#	n�=_Y�g!��E�����[��tB��Nv���G�^��;�ǱӊH�)$��7��(4��V�L$�l��M������6�N�LTrV�b*[�{5sPǜ���M2|�2�J�E��oJ�j�5AU�˿"]ǀMB� �Pة�@bK"�
K	�!XL�٦x�?������y��ϬC�I)���� eS�$Y��D�*�k��)f!?������͖T��Bdcg�1e�����B�C��-.*W��s��n`�nou,a�ƜǨ�q�0�D��{���b������{@��]���rE��fe���jrx�*��q^�B����I��G��Ͻiv�u����8w�V�O�t#�=��b�b�0��G�0��K�j.�u�����C�O𸿿�=k;���L[�������y��š t���Nx����A�:ؾw�������v�W�%����4H��7#W'H%��r�,7����.5m��<��;xyh2����@����V�!��z���v(�i��a~���8�˙R�P�r-nq����Q;�'��.hD$�V#��I�P�����&�5-�r��>hu{��p˜�0�sLwS��Ҋ�{H��.,G��7�[s�+�-��B^X�gf����d�<�/��S��F5�����U�;����u��'Rx�����E�F$sAD�ئ��e<���bTF+*�*z�&^�k|Ns}w[�A&;�/q;j�[��?yaW�(�?��3��͘�q�y���ޘ]��T��^��SP�X��,D8BR��4{dA孥��wBK=�m~�������b �pl���@4�V��*�x,�Y�Ko8EVP�h��PCfd���٫9�5�����n���}�1�k����]#�芻����B7=e��\���m�U���5��HH�>#� �7�����N��$4l�2z�����C�)����HO?���`憚]�����6V�7����^]�~���He�c��������C��EQ�e�)_�%��V�=��K4h4,��{�L���X�E4Ą���oʻ�w&ݎY!=b]'Od:C�� �"�����zI%*�X8)�a�;%5�N����/Q�X/����-�����=T
%Z��H�a����%���s�^k�9�C;όG�U�(j��y�Ųa��k�]Q�#����n���;�>'a]W���-�q���1�=�����܌'��5{ț��&8)��R��YL&�[/=��NQ�6]��'�$��\Asf�i}��'_L�v/��V(%��!8�(X�9��q������Tq3�n㶤�O�b:��љ6$%�y�@�5᜘�x��
/2���Bf78㛲�T"��[M{�������cL��o$�b�<tA߬��+e,����ۗe,��G�	(�4}Iz�F�ʎ�L��Kq�V��o��}�:�9�rM��o��nlK�J���n�>9]\xv܇����yE)ș��I�FŶ���9��}�%�C[ioϭQV��H#@�ȳT`�SBR�:è�ݙ�ܕ����������G,�Җ��$pgV��q���	k�S�c#�L��
��Ҫ�>/J�\Ԉ��oʗ��2o��O���>��?bG%�ו�܄�P{K���[�����ݽ'�ea�	��/���1C#�[���
�UH�L�����u�?_}X��Y�nB�q�8��ر�uY��~��O��?µ�R��w��X�L�P�ЛP��Cj�Jk�H��8P�'���4�ʦ?�ͰZ�	8���=�/��:Wڑ�>8m�aS7�l�3�� �q��'�ұ�߆�[��E���}��˥�ѻ�6w���=��S���Wk-�� �\�H�h �k��J�?�S6��x9]����P20\n��d�)�a�e�}�_S�����!��,�� j+=B����%����\}�9B�P��y�%�u4��ŀbf]Ts�]����Ʊ�N��d=���^hEO`�V�R�ou�w���w�EpQЇ��]����a�T>�&��n�{���!��jecE�����v3�##ԕ�5N:�P�Q��±<S��L` �7!�K�V1������n��d�LQ�Y8?�REW��>�⭃O��q��\4���G���ۭ���O�w�"�2�̃|U��\�<j"L���5�o����X��7�Q�xU;\2�ڰy��1�BV�Ƥ㖩�]T�1��?���Q
���(oE���;�H �S�Q-彮�E%A�����5����_k������ue#|c��5�(O���H��Ӵ\}�S\ܓ�H��덜�h\��s\aT�{�ن��$���\���c.��c���h=@�Asӿ|�(t��6%C��W
��_��J��a�	
�0�Ow�A4o'N��V�=zi���3��?��`nuJ�Mk�!g�Hs�Ð\Ώcs"0���o�'l��I�S��Ӆ�>��=3�����{��wf�������L�
׿�=pN��6¶ȘE`|�����e�Ww��T���n���tĮ��<�ư�/y�K��J7F����4�w4���;�Z�r���	�p�f'��E���T�����
$�釭y�D�&�;���KB�tW������}({��wiW�b��,�T ���A:��C�=Pr���i�_
E���vu�al���[��c�9����zy\�=t#��ۘ�5��ɹ�e�D��_�$*w��BvM!̟�����kzz�| �]���4��I3Aj���Q���{YJ���_�fdIFŀ 6o�����㴛2���^�R��b��ZV\q�:������X!m���n�n�x
���?u���ځ�Z�>u+�� �Պ��`���5'n�(-��,kɌ�sP��w��c�������gboVI*�u��������xK0�:�r)���<!rO�g7P�O��!	��Sd+��|55}C).���nZZ���{}E�!iL��+
���R�w�K���#l�	
.�ww��0��*s��<���	���Y̆8�ck��^2�X�B�&�G��� ?_¥R�x�r_!���?�z�!J�KZ��9��c:�qj�#&��X#�sik�� Y����k w�	�e�6��%��G-�VIF5�
K48Y��ʲ%��� ܎�g��"L�o�B6����k)�SWH9�r�Ǝ������l8a�;xC�hiM�����ca�ⷱa���Ʌ����<��S�+$A�{�txʰ\�_�a;���)�Ձ(6Pi�� �����YH'9b~y��ł���!���g��̫�]�j�j�4�y��dwap+��*����w�th��'�c�O���3a^r��(uR*�^�|&D�n��&�P]6-,�m��u�c6$ş�ǣSM�%/w�7(��cE︦�:�2Hh��U˛����[��aV�:�<5Ǵ��|j׺�edu��~{ z
� ����1�rՂ������L�f=h�_�q�v�����]��p��9}��ӒD}xc����	h]J��bz�4[���i_�����?�T��Eu��o�����xX��:�	�� mz	��]�/7��:����^��Ol�� ��a�+���	k.|;��m�F{A�s��t�P̥�yb�$�\͂��3#��b+�I�����x$%��`d�l�ZF��y!m��YJ3�y���vN�����I{r�0��ϙ8��BQ�~W�$i,���sM�ڶD���t��%)I�,���[DҺ��
�s����n����!t�o��awd� �NOu�e93�e���'��i�
R`�sOX��<)DĘo��·��c�|�s�u5�� �2:$#����膍�Ӝ���~��d�$�`����{�Ld���!�1`Pj�&�1����g������u�hr��_��eO d!�U�8J<G�) J��R�3�c���+� y9Z��f�H�SO�α1i�=k>���%���R���G~���z��)y���#'�����p�R��T��ԉ�0�'q¬������^2U�t�G�{���}
	�\Y?s��,s�����xN�"�[f,� +�h}�*߰�� )�g��#�w�
	zY�U�,u�-�;-�����j��D��@��R��Tq�l�2�9��י=T�ͨ��4֕08�(x��+�l x��E���b�,��ˌku�	!���?9��V�C����93�w�Ec!��r#�+#�ч|�S�/�Ɗ�ѓ��J��a�c�.�Nm�m���f.@+[���J��x���vy�תa#�i͚T�Oh�ƺ�2xMpD�y�շ��3z�7�w.��A��^V|�Q�a<�
[��,�8��.�4S6�A�XιHZ�|V|���qT~��{Z�w�%I��r��X佤I�zr�ݴ�oi�2c̇�t�ӄ��@���Q�'�㬾��/ �F�F��M�P�����Jf+�Xh+��&K�u�\��I�%Q{3#�0zl���<� k(�*�޵S0d�G�8�޵��+ W���N-�gpՅ��8N'}�4�$.\\2����N�B��FB��/5)��r6#���nu���ͺ�N�PQu�{(2[�Hn�:1/�Aj�h(`��	j ��^U��q��t�H�[�����OE����E�S��E�I#��L�&�p�ܑЋ!��M��~�V��d�ο:O�<w�/ �t��P�DHa}lq��kЦ1̇Bܙ�%x�
yk��k�1��X_��$���1�?"'m�Q�O	r;U����k3*-��ƛ�����+��-q����I�A�&�.z �K�~c�
�j'uۥ&px���:�?���s��Go:8� �{R;���� ��IG������z�cR_�R+�rWB^�hY�!L2A�.<��3en���2�����.Y�;.F�!�]wA��*��g����(���zB-�Yq�)��E������\��z��X�m=D�)�1R��ߚ��t~�5Xt�)��/D����D��S�>p��~��W����g[����'�y��`�~�EG���v���"�T�ٮ�l'�*���cpI�/"�0��@g��/��[���y�VyJC�M��-tH�����r񄭦n�̖�Y��Aj;�RyVs��Ac&	S��*]TG+I�_���ͭ=z]��6�y@DB�%?J�"_F*l�6W��I�z&�,Jodm)q��i�@	��>�2dE,�>;J0�?O/��ǽ|���=�f�}�Ok�2Lz��� :t��vq��^W+b_E)���H������cz�Q�<ũ�m�Q�iW�8o��'d�v��np�z�e ��e.�r���9M+����J�Ybr��O�	"2����[���+��).�(�����Pm��|��?1y�',��*��a�R���޷���٠�C^EӫqtC��k�Xhnwɇ��{�@����([j�dxh����vT_��AT�p�����L���Xr�+�H�:��P��\�Q/��ܕ������/��fA6�<�\�h��l�/��K�ey`q�|��4�Ǒ'�,�*�kF��6C���L%�'X��Iy����o�p�^�o�j�i�/||���gX��>�0�r	o��v�c�3�L}{�t ��H�X�=��L�}��1K�d���F�S�Ş�&�n��q���X)�XL�P�y��`5�	�������� 1ޝ^����������e�rؘ�ƥ�++�����u��pB{9��.�rB3Q��8�8���)]�%0�"�&��4d����v��SJ��E���� q����=ؑ�Rl]X0=�2�D �z��r-���ԩ���$�b/_�0�<�B����J"O_�"y���A+Û�*��ȑw�`&�����8h<@�󋵯*��$�E�v���E����\�b�;����@[�tJ��|��G}�'����u��")���Ae;����@��\\B��%�N(��f:{�'n��*�n�Ήg��=C�|1wO����|"7ml�#z�.����J�Td�`�Z!rC���X�c����~�W��7�/�z�����+�ir�G��άb#���iu�����P��$��=�R99��d~h�� òR��-�o��0rb���w�MٚD�W�"1th
	gx�p��%v�$ �r�,<Ю��s���ȁ��D�viK=uf�(���-���R�ŵ/'��	Rzi�z�G}%)��=���6��sSСЫ�t׊O}ī��HJ�=1{j���?������nc�F�����=�R�0���V#}�
�@
ep-t��-yØ��!�l`�6wMx�P��tU�[S �̒�Y����ɪ����x�w���Q.M�sdܦ�f��c+��?�Z^ȗE�u�ң�E�,S��%�N���<I����딿98�p5\���}��~P�󵧆A�ߕd��_���"�W�.��OC�喰��`��&8��e��e�+��͌�%9����tf��Մص�3��bm$�G [�S%'���z�B��Fc:qm�d�T�?oX�*��2"�}ϼ���}�Q��+���m��f��F���8,1#��)/XI����k}�7;��DYY�S�M�J��O~q>�^J��!�I�_�i�(��\2���*��V��	[���[�F
?��ɌP��f��>��+xQ��C�A�UY�I��7��١v�`��i �S:Z�DW5�-�����UnR�)
!��Ӹqӈ'g��,ô#�'�6������S���7�@���xeJ��nU���)\i��_�F�83��G/��8=���L��h2d�dQ`H{.��(��a�5O{.[/��R�n'7�|G�4L[d���܊�&!7��52b�u\�U��!M��"�~!�S�Μ2�}�)����.�+�\�%�]c �S_��6�����c�(��  TiO�T�"���:M�_�����p�b�H�|}�c�O�i��C����\��mW�U�I��:�F�9�f?��(����O8���"�wz�l��j���guoW����i�x����t5&���ӈW�1t�'��rǝ�	Ĩ�W���<;�T{Y����N���Ny�mg�8����ۣ�F�\�F�(�N�b�u��0o�!=���;�bb�:��o�6�ċm }�+�R*P��K`���G�~^�k���&:#?���t�e�i6iᵵ����o7�C3����7���Mr@�Ed\�%�ǥ��U�Tu�^'�^�&3� �2OW��	4�v��#_�����U�M������^)�#V��I�^��hj�K�,f'��������g�<_V�o�q�m헇�iL���dtq�Ցk��S5P�>��B�D���W�����%1��=�2ބ;q��ٷ^��yɸӉ���knO���W%/��Y��Z�"#f�
R�M�Z��ksץu�6�]��!�N�x�1���w`�>�b��"c�lۊasp�ݥD3�}�a}k29�s���-n�= �@i�3Zo�)<�,]^��氀�UWӏ$�fT��W�WvT� �	nj���i Fۻ!B�%tj�~��?�8T�)�_�R>bĂ�ʴ���e[��vQ��4��P��ɋ��:-)����=;���������w��G�d9f%�Sh����t��M�|�@��HEi���̕r�&�9�E���'�/�~�4ۼ����vY�i�.�"�]OQj��Ձ�;V�}f`Q�����%�HK;�^���-�������}���A.����E�i�?��4�Z�@"�������v֞iqk?��j�.s�]�Q�bc�g�v��N��e�I5΅6��5T�4��F��j��,p��íw+�ڄe$�ޕ�"�8=b�o3��G���ݚ���@B6�0_e(�+�w�����HP�iE��KԵ V���p~��84春�Ô���egc�|�S4�Z��C۱��6N6�����%(�3Ъ"�e�v�d�.�}Abt���A�|9�>#��g=6\I ��L��X7ZUzt��N�/R��C���d�[�CY��aoA�W��g�w���B�OHC���k���Z?[��7�Ƶsy.���P���ȣdL�($i�x--~�����O��z�1���
�H�`O֗Ш�.��F�����s��xyG����L�=Z?�K���$&����b�u�H�pz���/aF�LiK��g�c
f<xXy������y�ݞcb����.���K��!���.��S�y���iȜ�H;�	��k�f5Qp�Qg�E�	��A���׾,��<�M"���w_4L���8:�A�;�'R�{@�w�z�9�6�:�����^���=�G��)�Flc�����=��G9����}il��}���8�ٶ���|��;�U�CyzS���&0t��6�PZ���]]�T���:A+�{���72h���(P4'�,��-@6�Ӟ�����A�Z��I�?���)����PP�Ր��-	��%����Cq�vu��*е�3f7�6@�N#��Y�#U�1
����m#�W5����R ��8|lx���?p6p�B��-�S����
8��羘�ao:��ڃ؃�FL؟��Y��\L����?c,��|��%x�)�&�d�Vv�����4�IrA���?��B�C'��
A���>��b�z�/��Vkuj^�6�EK��Q�?y$�R�^�"Ъ��3��`���fB�[�6��j$U�/�%l�7M%uu "[����P��6�pGW���?���7wGC�pKJ�x�/���t�[Jp�!"dqyl�(s�&)�|-�&�f���Rd�G�*�&���;>�?ˬp�>?�=���N�?pw4�� �%���I�v�{l�AR�d��)��ܾ)��U��4��?���<�9^�Ƅ��<Y�Zk�<���H���v�/����~c�����R/#��*`��ЇM�݆EW��#@��o>���9ū�ٔ���M5]�	�_Ukui��x�5s&���Yd"�SfNp"�|Q��BD�xl�E��7!�F@��kf׋�5�3�^���$q4�E ¯����˫5(WdM�
�e�DMӤ�(�F
��?����GO�6>�X�Ș���)�ڛ3c
�c��M��N8ٚ���(imG��"!������<Z�{��%}@OPe٫���m9�$�%��M�<�X�)�K�x�e����V�ψ�2���v��d�W������S��
�|��Z�	�ɝ�H�ǞnwЖ����/n�M���|O=�WwPޯ!H��}A;+d���v"�%�h5��ДE�_���N�YEoe�WX��a����N7��Fx�T�F�6/�x�&#��`�����ra�=��g6�sI٠�!V}=,���~�Yf�j�i����ݔ̜�K�� ���ں4p}S&tql��fI����Q����+G��v���|�1��8��3�ǋoB5�G`'��ghAc1��Xk��j>���7�lJ��eߺ��%\�� o�_�-�R6F�dW-HlF��?���-�?X�:;�h��s�Ȭ�Z�=�'`�,S$B���ˢHŤ �ڢ�?�IX��DW6Z� �|�q��{���_<4d�����������)�I�_:N6��x���Zg�'dcNH���f7e��7��?��_�dbl}3���D��膚J1��sVJ�c��wz�����	�����lV���P�^�ں��/:� S���ʹQ���sp՛x��:&L����Ъ��;ӕ��a~�` ��|L	!S�Q2V�S���k�O�W�w�QtC��C��}n���Ȃ���D�݉:������s@�^��~�)���2�A �dHCj����{��d��n�%�%,���ʽ�#��+�IG����?���jǓZ��g��k��n�ʒ�.��|Y���8v���}���	X�j&& F���q�W�!��p��� �x���|L�'T�"�0z��B6�Q�v��-	�Ѡ$/��\cU�k�E�i}��$�ݗM"���¨kFX�R8S����5ə퉥�<���/�n�~v��&��Lt[��o³���x�����,T���XG��xvO��aP�E���'nLE�W��D�X�]��`�)\D�Q���Ř�����׵����s��D���|��L��S�L���n�DpG�I���e��c�����cU��N2F��ZN�3���X�����Ց�"
�4�V5�Jf���6`�����
�BV�'��ݗ��C7o�\�9��wZq���[�+CY*y/�H)1���V��H�;�8n~T4%�&��K���z�j�`���t�e��`j;���q��#��j�V%0�����.�+�ߟ���0�M4-��(�����s�����^�2[��͋�J��$'��̭Ƨ��`����'T�n�OB䐐�/��\<sۯ�#]5j[$v;+���̷o����1��GZ���rI����t_�;J���z��Д\|���G��ƢF	�t����S9pVfp����tҞ/u�W� Fx�p�J=���!�<�"!<d~y��}z�u��?�oTb�!(����}8��)g{��@'������T���W^�� �Y٣.]I�@�����)6Q�O��� f}^9p}�O�	sla�=�5C �0�2��F��e�ܙIʔ�)�O1}��
�&��g�w�yf�&Y����o��[�+z�����t&��\� �J�o4�=q�!�������؂��̳�����Ҵ������SO�5}�# XN�:���Aj)�i���I%x�eL��D3S��C�<�Ŕ��ͳ-#r\ts\s��������|P���\֫&7�o�r�}
�]��1	����x����W�u��=08)��h�=�@58T�{�ֿ��a���/^6H�I����	�^�L�O�j��5��2k��Dz �WL�}��3D�!}��p�Rx��N���O7�a|˰�y��Я+-8Y��g<7��w?��/��j�;�#e.V�R�R4�3m'�x\y��Yf����ݚF#�ڧ¿lAsD�!�_Ϩ�A�̖0e�@�#=�bVrW"��x���*��M��.$YEz-���
��Y�IY���1[<�g�L(a$��J�ψ�5�螋cY{�jU��S�&sX�n0Uz��������A�Ǭ���OEt/�Q8CSD���\+�p��W�S(i<��<��U�-�Z:Y��]�Ht[��%����1ŏj���$Nč;ك����?k����!��.1���
JDc�"~���.���ɀq:��սO���}	*n�q�L�l�P1�]�����n;�$�4#z�c�M��yb��,�8/�������`C8@���f<�M�6�hg�a- �	�nL��y`֒�@M hf��h�}:�.��;�O���L[�W���$<��)CQ.=�C�zG"��dV�=l{��uu��HI�ݛ�Ξ�Ե#t;c~����"��SԇJ���{���s#�TQO= �XE�~���!��VV�Ը���ıkE^�0�����xh�)<�h҆�X̷�}il��@�x��d^(�1����)��+�n$�%�v[?x�J�J��: ��ra��o߾Y���t�{�����&/���X,�^ֺ�I��Æ�K�7�v+NS�t�XXqG�����?�`h�HW��$*�����h8�{ ��l�_wr�s��v�n��dz6Zi�Q��/�����pΩ���t<Wr��D���(�Ћbm|��-'!֣���y����ߴ8C�e��/k^���P�F���6ޭ0���vɑ_f}N.ǽ����w 1KX���f�<L��R�b���hcY ��|���%[������	�I�.~`�A n�#;�^�<?�<���X��>��G���>�F���p�Ɔ�o�!������W�z��um����[�	���owZ��i18�@�uq�W�S6
`*��9�^��� 4�ZJ1�Cy��N�����Lf>2��%����K�"��^�����&dO�^�s\d��\�8��wX���8�i	����U��W"I6- �Jn^���s���Xd0	[mp���a���F���,.�r�
���m��z@�`���v��_l�b�ӱu�ce?T��m��>�̣�f�jډR�K�T%bS-���A���3آ����<��D��S��\���/eD���_ف�b�ax`d�1�{�.%p��[�#R��]�B�������Y��Wh��#�ʆoFS��Fi��zc>f��L�ΐ �B��]6�������,g�$"y��KoPR���Ť9��8@��N$�d��u��˳�c��1qsz@y�Gb�0O~O��%�����=��b|�<!sznEX6�kO�J���Z4�У	�҃��X�?��?G��b.Zu�.��$6�1��0C���N�{1�Ύ�7w��2�52|���zQ�g�!A���)���5�!��w����c��)�q�
��	�K�o�7�X��0��8�8�!v�4�����q�Eþ(�pK��#�����B&���{3-��C��"ȶ�[� Ѝߞ�=�}娰�Ăa���jԚ����
z�yv5l��;�G��hA��g�"��tq�P��VRM��ƻ�I4M�
�����".���m��,
���&�GZ��ɒݲ(O��R��R��PЌ��C<�ͣS�#�OY2=	�Ϫ�����;)��.g$Q���{|�� N���ʹ{z~'D����U���ca�[�m�w��`I��M߯����!d Wf+넍�4k�Qej����'�?��aZ&�,�ش��f�����Nc����T;Qƅű϶\����/�D�+�B���YOH!�L�����3p�h3!��G:�ܩ�w�k��JG Tyc������~�+c�Ѐ�dU~�c����fq��~	x��z�ߧ�NI�P��|>��v�a�^��"�
{d�2��RK��W7����$=�t(�/eWOGj}a�I��-��_��QWZ�U�Ȉ�:
IF�t ��R�}�5Ņ�[r���n³m��i�W�\���>v�Tf�62Mh�T(+��`k���j�S �/Юjݔ���)jQ�!�HYFiA�d���i��i��|QU��X����-�<lkU�~.6��q���î����ʎ��:)�°�)�i�����j?�ѷI�� 7���V�8�]�t��]<��º������|�Y���N��2/�r��:U���DJʶd}�KyX̖�9�'����R���"ǦEf�Qǿe�wb�� Wk�,�G�5�`�����3:E Q�*���Syv�@��CD�1����]��$���0�_�cK�C߈q�ui#�wq�B��Ώ�V���������4��E���B͈��#��֤5d�Ӝ��r��ѡ#U����r ��;��^�ͱ�w��k���1T�X���|wco[[p������U��=M�#gt(Ǌ�\��f�R��eY~�
!��=�/�dB"��^�T���,�z��]� {36Y�Foo/T$4�%
YÚ�Yʵ�,�����6�ɝ�e��.��Ʃв�[=�8�������}��a�c�P�\2uO���vܷu �/P1��]��V��Ե�����3�#7n�����ߐnE6���c�(F���BӢ{ѓ��F?+K��6���]xY�7b:Y;B�6u,-���r�$���:�ʢL�˖U0ڝ�Jg�=j��>�E���6��֠��c9�dx\��k���Q�4S|{���}�uه���-u� ���%L���'������U�&���=��B:�ݠֹ[Z�w���Q���b��S:A,/*��t�fwNrģ�&�8�u[k\x<��@�a"c���B+5;��#��P��|e���!
�*��t���
�
�FT�^V�ǋ�S������a�(�֎�O��q>��.���i׭�U�R�ƑqE1����i�}������=п����K��7*e۳X�i��5[���ud�0�;d��׻�b�C�]B{�2�}Y,���%�.�e:�;i4�v��ʐͮS�	~"�2�|)�VX]������a���ҡѯ0���={�#�v�]e��Ŭ��oS~�,H��D6���j�$V�\��IPiX�ˮ �2��+����.�)Y��:����UlǳJ-ӽ��Y{Tp��ʅ��|?�_���qO���@�'J�mK�=�~MxB?�䴭���@O)m8�ۦ��Za-���;�kE-2�����d-�č����d����[�\��=<�-����'��pe�T�䒣�9�`���nV!n�1�Nv5�ʃ_���P5�Y�2ƻ�X��P�6D7�HY��s���Ր`��4��F92�˕�Cҡ�8`��� �5�o��
$�Q�Hps���?*\7|�Ā��+���z[��2��Q�!��,ޢ���m�$Y�-Q�����g����U�O����@^Wl؃�jo�������R]xr<�`*̘�P��#W���v�������A5����ɏ��]�3<b�f��Q��zP�z���D�Z�E�?�g&��2��AOߠ]�k���9?!��d��#�D�a��<���τ��gR�ˢ�3 ��?�2Fy;��}����Qf��y*����s~�15��Z��G�$��x�5�T_��\6���s�W{��N�d���HezL���k��8��皸���Kd{�^���ٜk��q�F���w7�}ٳ��m	�m�2�*�[��K���Kܱ�uJ���~�.zN'���Y$g��PΊ�-�Z�����F9}v-4b��h�s�������L��Y�N���!@Br�y_k?/ ��0�D�u:�w��:`�>���Ԣ"��l�"E��\���o�9����L��]Q$֩跏�郟�5O��S|�/���$D8�2(D�h�7>sM�ϭu�F�|�>���~��"�����RI����Ӷ�XUx<F�!���V��	�iCfdE�f�e�P�����:��������^�뿓� �V��3<�����cg��ˮ�F�Y�w�{I�a7�a�e����	r�/zQ�+$�3?���~���Z��P�>_�-~6�j���h���|�z����4�z�yV#�<K��F6�M���.���X�t��p�hV�]*{�%LB���H_��.T`9�����#�zɓ��B#�?郦�������S� <�CEwbQ"<�R��(S�H5닄Z堍N:��t�&/�d�Z�;�wS�?�ZN}��F�FS�nK_�ج, ������_B�&Ƨ3����?���j�=�7@�w��C���������Z�U3{Ow���1Rʅ����[�.Yj�g���J�)�[q�@
�j�-��[xg��?�!��qn0�^"�d�qj��W�EW$)<?	��d���*�3f�;� f�cҀ�un��2�� ��"���#�|G�����u�_OAj���mUʪ�g_�X�I��MLu��u@[}N	'v[Ui�&K9���-����٘�f6�?��R�ۂ9O��ġ�;�)b0�B,�Y�O�?�YV�6�`�[%�o�y��1���)�	������Z��DL�Ǎ�zJ	M��w��|U�������#a��C���^,%lc_O35V��;�%��Nb4��Y����Ketɛ[yVP�V�-�k�����R� �׃���ÿLؑ	��bU���t��N�+�#`R��	~�T���{���:ݹ[�b~����0x�P��&�x���s�@�GL)j�'�
�����
���i� ��cΆ�w�$���*�B�#� ]oH2+�&������{���>���b)�_���z�5,4R&��M��u��dY����(`0��Q����#�5Z��ú������,��)}�b\M�)�|L�C5��%y�.^�����Or��F�WW�}� � V"�iڐ4K�rd�����G���T����QM�Da�\�  �w�ԚnR2;�O,-�+Ȫ�^��.ŋ��U\�͠3��@"����? ��Y��%�N\[��d�
��%���\S��g�b���@���a��f�i;x݂���Z�NU�5}�0�҉�]�����S�U_d8��z�v�Ԗ(.K�V��T���C�6>�b�S(d��r"I�n6:l���o:``�ﳽ`���ɐ.�IR�4 �%��P
���yV�g91��f^�Ƀ'#�MuH��$9���v��!��Mu����i3�\%�&_��"�l��3g�a��IB��f�ToR�-����G����7�3��� �Y8a) �9�.�(x�M��@}Z�m��mOr���u��j׈��|��2|4XJz:K\r�� � 8|lTӧ���9��	����[%
�ou���1�K�9k^�����w�U.���<��ee�)K�,5%��2��L�ªOd���Dk�����)7d�2V�;�C���no>��!�}҆��/���h�`���� �����s/��#|�-�����ݖ�w�MGE�7�������gƲfY���
�����tG��T�Q�=�= l�zl,����(�$��P���4��.����^���8�6�o�7
L3��f�zZ�V����u:���œ��.��$�G<a!CͶ���|M�|�Sr��g�'�*M�<4D���������A�^�B��$�f��|�3��M�x�"+ۓ�k��BbS+\�+���E͛��1ժv<�ˑ`&`KJDLHp�}F;�|��a-�
��0��y�VQ��\k�z�=�IP�]Ni|0��ÕR) ��6m4��^Į*>���/� W�⒓�~�&�t浶R����r�jY��jD1�M��Zl�\��H���,둱|�`�nt���qP2ق��0!��;���%�>V��(����ջ
1S�G�����v�F����1��k G>�zl'*�N�����ҝWl�v�����"emZ��ڀU�}&!S�����#ꑒ����.��=�}^���$T��
��|g=o"~��/�b�g�T�J���I
iX\��I;��D�CJ�(/9�b �S��|&�_�ҽF*o�-������+M�S:`�V(�욏�Ĉ�̿-��KY�V0�}-	^!���Q�@��(�pk����țٻw0� ���=�������'ȃ��P�ܙ�|U�9��30;��!�20l�NH}Q�]�S�2�pa
���V^��3��`5��e��@����f�k
X�y���F�y���hv�:�vJK���S�W�K��ݘ��WC�/A�@c����y�@�¢ߐ!��l:��]�ᰙ�)�S���S�3��}����Ĩ߳�CY;5r	��a�4<��P�B��3T�ȟ�n����+�
�3�>���Ȋ2iSH��ޚ诖��Q)�5���u�SM���2������Jչ�&pb�Œ�;�����m���_���G�8�)}0���> �"��q��!�m���x{��Ƚ/f8���߆���I4�/ޭ�����&�������i��3S�6���
�"��+$��R �P�`�$��i�\)���UN+�
�������.+�7�5������59��s���I�sSu����e��H��u-���
̶�<����+���;-��~���"��²FP�h�{@�k�T�W)Pp\�JAL�^��&�Kri�_
Y-x��Bc��7l|��2�-"��Gg8g��{��n�G|�U㙤�$�@7�l�?�Nm`(xpr�l�B�')>�A��pP�@
{Z/���KM��n��p�J��A@� v�b�J���a�X?�yJE�Y�d\�!��m	��¯�Q�aEY�s�C�K�9�W��%��X�gM�:�����i����}�2����_ϗ�z!���9��ܛ�I��>^2(��П�U\(����i3�6��;�	���y�ūHR����]�"�{���������_Vh[�sJ"w��-��������Jq�p�V�֍l�=<��Q0�a�ڙ�0U�{d?ہ�?w]��-�U����By#2�r�ۜ�uXn�N=�M�a��J8�m�=�6���!�d̠�����^��\1F\��-��Xb>�B�X�r������2��e�s�	���!��!�$X�G��,]{@�l1��~OD��C��X"8�P('dS/���h�����CfM��1ΛM!�J����-g�>jOjn�'�⃻ǳSA����w����*������@�^�u��f�ϫ�HE���i�!kiʤ���Pv���-$Q�<Ѕz�fW����vF��%�t�������]�C�;���8`��ML�iYs�v|n�4��1���⽣튜Ğ���_�>E�Q�/�˔& �QJ.��!�k&�<�#u�TjPA]�/���̟I���u�^0i}2E|9 ��p�9h52�����c)��r!��N�$����V�E�S]��ϵ&��XΩ��[������M�h��s"t�K����w��T���_����tY-����bV�=]���L��h�K2�7L��R�Y5�U͜Ι��Θ5�s���{c�sc`}�P��jSTH�(�K�X�vE*�r�����琬?�=��pܴ��� V�6.�7=Qt�ˀ��xf1��r`��gve��7�Bv�*�F�_*����Oi_�}A��	}�������Q�Z�/�5 ���Փ�ڌ1?yf��(�;@�>����"�ӿ�Q��a��D���0Mn�j'Lgs�������bo;D�-�'x7"bx���?�T\�#�)�X5<��B�������R��T�KZ�h��������F�Y�6� (��E������W�i~���Q���y~J�S�◼;�#�h�!�͋x�l;��f>.Z��ٻ�Id����ƸF��xZ	��U��bI��F�'ա����w�e9�V,�
;4���U��K[a��$Gy}xVk#�y���_qP|kc�\�٢��-��h���a35#����1���o�M=̉ת�]I�$�?����1A�������Ѫ����z���%�V��S��:����Y�	U�b�c��}m�7H:6?���4$�^��2F��n��a�Aa��M�'�f9� ra�}��e��jC��׊�	U�0�H���Lo���R���"q�7�P#f�=���J挤��`�kx�r���y	��f*�*
;Z�2�	� ��|LZ��B3һ�N
��=�˅ �.Q���5��ĩ�3碭c�]��Y�RbK3ݤ���е�~z�PM�f���7H2�ſ֗��޿Sb��K�4���O9V{E�5�5��@P���O���I�e�#��� 	˞��xw��0$�v���y/��(Va�7+����v=e�ÖљV������P�s��ҵ�5�#�>|�˰� $O��6��@�K�@:�������O#jgE�����^�4F�h��*��#��� ͿZ9�8(c���zu�r�k�)M�Q��^5ʜi� zС����:�Zצ�E�)r�q�����c�/^H�٤c�����d�K������4В���ݧ	IcwD޹! �H��i4_�o�5$��T�;�-3ց��?-�\�������jGv::�0����;��P����_O����0i�/���=z�"��Hi�o�����t��7sBh�D�4ݸ��!Gi�3=�+�
k���{}�L^���{h"*�tB��߿߹��L��$.p���tU�J��<��~g��~X���#���9n��{B��D�/G�V�_��s/|�=w�*�?��B:�N�#_|��FXGX
��E� �#�b�.�{���������,���XP�p�ߞ�D�}f����NqP����[��`Ӧx�uu����P9bD��HxvǮ���,�G^������|�Qۅ@hKi���L���Q͠�U���$��l���r�#ǩQ[c�0>�9�ϿQ����m"
��%xc�ˈ�H�I:�n�ϵ�5���{f�g��M������m�cϸ�Mb�N���*����V WY�J�f�d5�t�G��J({aPG�'i ��|-醯`�ϣ�v�H���Q@���BK+�қ�2�γ����Y��?�@��y0�-*�����*��.o�H����9�r��4��u�|��[�����H���:DG��i]�*[��>ٺd���$]=�oΛ���+
$��sq>\<�5p����+�> z�a�WC�>6B��#Y �A(���-���|P�jI��@�P
P*I�ː�������h�2O����������-wy��4�U��~ֽeG��Δ�#�+�w���R+���+�N���PJ�J@�����0�r�g"?����d�:}z���H�O�]�-�*;�� ����NP��tݺs�V���{R���ZV���MG�+���kM����c����Im��̔��+�	_C��6ă�p~}i�[�B2��dZ���n���F�-�/5�%��=��ѱ(�����K�z�BQ��@��@"�ˣ�~�5]z&�+��^җ=��VNsty�^�$�&9�k�@��u�\p�e�Tn0�%�Nnb�����Q��������*����f���=���H��ZE�"��oS��
�0��W�A-	�ha_#�UF
���o�P����r �($*�3&R�`bZ��ν0�C|����V�׊�L�F��Q��3��G(3���<-�
�` W���o�e�����W����S/�	Q���"Ϣ��ǎʵ��:��'$U�����1�e$��@8����	(�lŷ��]��z�쨎}��8 %6� �S�	Ae�74]��Rq:WP�:-�fb]}YL�YKcsN�EC�X����(yv��2��9-Nw>� /�w�w�E�Ýr֍��Q������v����3m�zx��*�H
Q�Fx��6f�~[y�����<Ә��GBz�V� ����2;ȸ��G\�����N$��Ρ�-)P��X�ܻ���h�mq �wz���D�7�q��2
���pt�oPj��1�u�bB�8��zu�:41���mx�_��B�s�(��zgX3L#Ѓ��"z~.F�ֵT�G�fǺ��<�QKG@�C&$3���lW&|ʥ���=]%e�L�撑���cwg�3���f���$KC��1�m��$D��,2��W�t<w̋�J��Sw�J5?��#� ��Z*�UXZ����]��'�8����_]�@m�$1�Bi��H���;ψt�\�q.���HLċ�FJ�e�k�%zߟv�x(*��s��x�r陉�~.�'�Pݺ�$P�Bw����\yD/�m����b~D"�\�E���pV����:)�$N��e�RjS��Z����0�B��o<*��ʊ4H7��<=�@�պT��j=���.��vt�T3& I�}:���?�9�_�ќ�ßB��@y�n�B��f�7*��5K�Ṋ�$�?'_m_ߐ}q�2�h���/�@0�Q��:,���|n����.D���tlN�҂W<㠊���puc����N'k�4J��D�3u� /@�ɆE�A�ȋoO��K�'v���02"t۟� ti�՗�1�&�`�2���`���r�KH��#Q+��[zrzBUg�%�;O5��JM�I�2�8��N�Uۯ�<��g�˶꓀��4��;hJ4��؛���ʛ�sP;�.f3����~�Ѱ��_%��dG�틮;�����u�e�|��]�p�DwiS9�4xh�f`f}=,V!�ܟ�'�9D�:�愸J9+-o{q�u��S	�H�������8�M"��vv����1v�I������@�#~�))cѨ�e1F����:����0< ��!�E��rZpF5oQ�djE������?d`o�c'�c����E���K���a	y���1���j�L�m���f�Q$Ϥ6�aQB���<�e��{aX
?f	�C�L;�~b�I{փ���5_�\s3���(;s����NI��ryg�v+�:t�FIX����}��_��}�<�cOY�"o+�e�ݥ�
)?�!��*��[��v��Ţ*���5L�����CIgv�v�5p}�s|͛l>�W��ԲP�3��}���tTnp}#�^�9�[�Zd��	�����U'���I:T�&����=�u ?� 9��ꑝ���g��
g��:�S�!����y�B�f��Q�2/�}��4 �^N��z.��iz��CN��d�1#W����۪n)�p^�+f6c�S����/g)������/�������=��*���f1�־�$ ��L�&ΰ��W��3�)��;pf�m2p���_��B7�o�ԭR�EiTՎ��,IVH�.�'��B#��W�Uݺ�*�C����~�4�n�r���2�JGy�"��{�V�(��d¿;\�i��(&io�%��?�����)�	Y�:`��7�Y�JW@���t��M֬���ȏ��S"�(r]�4��־=��.J��ݬU�X1�(84Y�)�
���:�}-@GZx�������d�>^0�ZB�W�q��7E����Xu�]��d*\�6�+�ْ��� �{�U�l�|]);��_Rj>��ncQ�Bo_
>�8v��hAql;9M�s���p�%N-�#���F�)��j��Lm�ߞ+*3��\�y��ƌ1��\��TZ���o4�AZ��w�rtXcZ�ɐQ��S�>�lO�T�l��i��E57*v����Bdq�<�����#>{w-�<k�>J�g�|~ճ��BpAm5w����Iq𯎶yg�JN���j;d+��;���ƨ�2��%�vU���l�^t�b��s?�O�ױ^��->'�|5o�D�&�Sly��w[Y)A�O6@ӈ�\;p�4AB#͟�
���p���.)g���A��[�
����Z�����ˋ��� 9@����C#��j�?�a�t��.ܩ��S�c^=ï�clm0���{��Z�ki~a̮����i�J|L��3�ʮ��@b�G�x�]v��Y�*�΢��uIC+{��e��'MA��wE'�)q�ܖCd�4���i�/���'WDs�up�P�p]�O���q�7 ��@z�vrh��ݵ��w"�]|�q����4CH�`���aE��˗�Ymv�~W+����Q�b�+��mTsJWk\g�;��G�'��e���elo�o�a�vf;\L�` 1�&$��|g���?X�>u�w�sôxa���f+xz�L8��*��uԲM�h�%j\�Ӻ��_n��3He����i�������h�B��61��v�N�p�Oj\�(���i"m�i�C*Cs���� 9Ǌ�t���œ`u� ����bb�V�}#�0���1s��oo���p��>|[g$�[���i���7��,���Q�D�L8�X�/���eD�鮼yW~�"�>~�ʸ(����gR�P��!G����u�<����МM��F����$dlY!��~N=u���w�C��"�pd����0׿�(���0����7�<ŕ�����ڰ&E	c�9�C-$�?��'�!)��M��v��F�)�N�Ϊ.�'�΁������l�~�x��Ս��_me�cU�7���./�3g9�C�P����q6n�3W~��b!�{L����VJ����}�d�ܡWj��+���!�x���+d5�&����&R�|�t���*0����.O�Կ^���~���3�X�E�r�U,~E� �j��J@��X���!�m���;A�n�� ��H���;��]�2e&���L22�k�����,��Ó�3����,���c���s��X�h+�fL����+�;=��}�#y��;*%Ō�ڭ_���AE�J�-���0d�ܔA�I�걷��l��K���x���������^ò�4�V���5c	M�������6���^�B>� �B
E�Ez��-�T*yX.9,���$� њq��ݾ]	������>�d���gX�6 IB��m�#K�~_�P7����j����?*�s��C;�CWx����2�@+��\��V܃��+�fu?���@����{a���ä=�)�6��k�;CnS'pĜ�� �5a��v��
X�(�����:ʧ������+�X�鿦����:���w
ţ�Ij֘3�"*��Z|ݓ�/��a� �L��4� qZ���Ѿ�!�tiuM��`V�CB���eM��I7qv-�Tcg�TA�88���胶=�H
jć�"���3IVG�y��jg��t�kR3hI�ʼ�$���>�Qz�2sU�0]s�5�_�g}Jl��xa;�w�w/� V��#�k��WD]�@�7P]ߛ0 tvj\�r��.P*�����m|���u�� (�>E2XI�\B�R!�9��AAЁ$4ǽuA
�J3��+�_8ş%��IT�y��H�5֪b�y`��IE�l�D3�f�O4)
�x_[������]��ѭ��b5�󉭍��Y�~E��F���>�缕|�A!���kwfeg�}�h�3�K~A�&d'��QBe�V�.՚�<&�]��|�#=bc���t���+�+�p*�&���Prw�����|����L\S����2�}	�(���$��$Z�F�,�Nth�^�m�%B��k�QP���ǁ`܎Z��je��G��=Z�|)�&�tM�|M�舖��u����tW�h�.YL01_z���X�ww[���C�C�h��:W$�R������h�{�?L\h@O�N]�U'�W�̯{���3��b�X��b��\��K�_��G�@�Vk Av��`�&�6JE��B�n� �g�M��]�C��y��<2֞����ť5�G�������E�^/�M�Q/���q0�<�۬<v)�W�F��Π� ��J�2�6��/ʲ�+?���x�x�* 3�<ϤJ����n���U{�2Jo]���2�.���PŲ'�D��Ϟ�X3�`��8�AWD�_̢x��-μ7�����b�F$�@	�
0>Z^Tvǈ1������5 q���C|�b���0��� T�ZgFSo��v�xB���.���A�.��Ec!���|���7J��֎���%;X��	���ey�$a�[	 ܢB^<[��uc"T�ca\�`U7�P�_�՘�2�<}��΀LW�%��R���d~+m ��m0��B�wJ?x*��Pf���|� ��E��b��Z�^�{B+���v�h�&_�^�Fi¼I�Qt�sth����&��=q�P�O��q���*@��Hl�>7rVJy�ҞҰo�/��Q��uy{�y�±H^6)�"!����CD;��Ϸ��ݱj�pE�hQ���dp�!�B�lCq)Ĺ��7c�wx�/�otH�����M�UƝ��nT:��Z�d*����	R��}�8RE�Ft���|M��w`�۬E�&�f~���%������7�'�ݩ��c��\�k�����Q$]�Q�˭�X�ۺVK���{�l�ܖ2��J�<�mGW��]�>����M\[��_�fE�Q;n�Ƀ��p�d����F�tx������Iͧ��4�:&e��'�|A�H��q^����)c�)���M}�q���6��j���c�:��2-X�KcV�
�$I�j6�=R���T۩v�V�D���K�~��P�J3:U����^�%���P�yI5��R�}�/�)8�����/�z�+K
rQb�Vg�ҭ� \2bMNϴ�E��]1�3Цz~c�XS Y�����ރ���R/��2^͠�߸��Z����>'�
�!wLE yj6�?�����o�ƶ�.r�Bu�	|D3֘�?�MF�	j����Q2�Gdn�[%�|�Q[} �	�麱�-�8;_ە�-��T5�=��
�h�3�I��b�_�6p�t����|�O<D�3E�=Կ�M<���5�~���y#C�EZnr�MpD��ZM��Ҕ���[-.��"��[ 8ʅ��݄R+�������1u����n-�%_�d���X�,jn<)/hr��(| Xib;J�� dU+�n������U�W�ԟ?;XFB<�Z�4�b��nn6����3޷�¤ioܣ?���kRu�ë,e���̘P�n�	{ɦJs�'40<A�E��	�L�l�������M��]�U�ڪ�����kO�^�)��փp��W[�7��. /	3�������$����Zn��
�[�^���Ay�E�����s�"����E|7)Q����Z���l�k���1��ەC��d�.֝���O���-r��T�h^㗠�~�߰�C�"X���A�R�S�x9�q�;!��f�~��-A~��YǶ��jP�I��l�Ψ����N@�1�Ə����,�¦Ű��J�g8�9�_I���-JM
��'6��4J�Z�B�t��m��O���M8 ?L����$[Xe�7�C*1���6�T���ŧ�4�N@Z��m��ˀ�Q��[=(��d�0�ɨ�]A�%��I��>x�J��N�3`�9>	B����6CXR��f(��~'>`#�f؍���n�En��8=�����{�F��.�Z��[�3&4�B�:�!�������~9��!�E��(No����ck+�7�9/pm'��Sv�b�����b�ЩE��a��K�Q�ö4��q[�яJ�d�#�Ԛ1<rxh0	�+.�Ԕ��;� ǵ��:��OH��o �u��.��İ+u~�6d��e��q�|@ŵ8�<3R�͖�h�-�'��t�T��M]������4�;6�6�r\�7s�Z�]rE��U���7��Oc�/�$w�f�A}�+	S�PKK߁%�i��^���d��G�(Z.�B[���N�[N@�H�/�����]�qr�I��!�H�+��[�����Z��\Z���i�hv���rn��J��Ԗ�~
�Z�δ�ъ��ݤ��ր?U?���F:�.���y��?�\n�+��3?c��!L�Ca8��S0�}	�I�-�P$�dxV��MMD� �EB��?{� �LQ	"��,����5�urN���'VC�{��L��V�/�K�uZ�
ҵ�xm+��X	�	Ov�_a�T��������T3�1�~��z#�gH�>�k{9�B�DHj�DF�~1��G�6�g�C	�Ϫ��1������I[�M�J������)幕4ۏ��|%ʯ'��ǌ0�^�l�: S�rO�#!jW��.�lDe�\&2N�Њ9�۩���hF0�u���!�x\:��y-�&YJ^u���{�����z��$�VEs~9���CO�ͭoj/㹚�=��[�l|:��C����9 QO���F�{g^���I���P��|�)�t�/�G���ɨr-N��?Fz5]Cs7�1�����l��s�wk�#,�����r����1n�TZ���7�r��H�>g�g�9�ܠ�=��#X�Y�ᜍq�*$�@>e�7�u�����a(�!����d�/h-���;�?@T����e.%ӊJNm�@�-bF��&m��amu�\��n�n���/�� ��c�(JwD죬7d�.���)3�MV�!���X����u�[�c�zB>`�+�6v�v�`�팵�x~�\2�����»0�w�I��kڭ��+��'q��A�C�B���iF���]����(���Rc�o:��/N�+2	qNAc�=����,��)&��)�oȏ��P�
�m�9y�1�(�����X��~Ӫ��UhERϪ���x�	鄉�/3��_x�z��82@`SJgSO���*lWQ��T�8.vۮ�uC�pz��i�����6���8k�4�	�Lf�ݝSh����U��(�)pA#�B������r?>Q�G�7�Cm4v_&�z܄��
�50Ÿ���s/�q�
&�$Z�(6��2��fZ�5�|8K��J��Ȍ{d�/s�ErP�kJ2F�༽ I���B��Ǻ;�˗�Ñ�i+K���d�_�Q�Bw��1n��r�8p��8U�	�ֱ̡@����g�E��6tUp48�u���`]m*ߚU��&� s혔C7SViD��ӯ�х�<�����|Sحe9���i����2�{W�v�p;t�'Ҿ�!'�A��s�[�0���R��z���γh�9��[NF@�4g�*nK���ci'e���"rCG�����YC���H.�T]�n"�B=�3�5�;���ў��TP')<s�Me�H�����b�, fr�e��O�٦����;+�nq+GܡS���"G�>a��a�}�LN7P�C_|����-Ef���)9v7�hA��$K�j��d`���,p0��S	��݈Ğf�o�����͔��g�:��t��|�(ؕ�����6����._Ѽ�b����#'�i��բ�驋�"{�K*��v��_�X{�XBД湥t��nq�ڋ�M����/XA� �T�jR	�c��$=�����v�_���,��y.����~���v3��a9�3�#�Q鎵d��=�=���M�E*1��n�nK�Z�~g�N�R���a� ��$��OX2�#��N�n*�����?E
�$����>BY���TB�m&�`��k�x��eV_��v:V��
O�z�gI��cѶ��`��*I2��G��︕�q��M�Yɻ�a+��X&�p*<U��')�N�_�o�H_XK���jStU
 	��G�(��P�H��=����_��1޳m�f/�G����)�p�}'.+�oP/(^g�o^)|R�El����'A�_n��2�$��/3�E�a�6�,@��d�8�KwF ��.�5ךe�\�(�/5�W��H=���	�,������c>o��V$���U��������5�\��{`�+���g�W~s�:�����ɝ��9V[�|�)m�ux��-���
2q�ly�._�Z�XP����������:��n�,ӣ����]�3�Q���
�Y��UY}E�ܐ�/L>�(J�al2\����bE��������! ��0���b�ޘ���R\�`�F1m-���DEa�׹Й�� �G�1�weE2_���n��$�8g�e�Pż�qY/ҷVq�O N�����MZa��'��#4>i���҄�3J�=4��I�, �kJؗ�F`�7��.��j��)7ָ��AP�3�I> �br~�7q¹�C�Ǻ�����k�^?<X��HM ffH3YH�3���>�`�W����߆ލR����y�E�4C�J汨c0��ְrp!H+�ϝ�{y��Mn�:��e �N�*&AΎ��'�͠7яO�}Э�n�.H6~�y	{��NJ�Na���sRf2R�7C��c8�߉��"�г���)$��@�7Ii"˶N�^^�qTZU��d*���+����	:A������4]�Kf�Tco�QvAѲB�v A���.��P�Yuï�I�����S���H���^�iK�9��Er�݅�D)�!�D��(a�P/v��V�����a��e��Hv�G�"A$xY��$
܅�m��*�@a{ML*S2)L�ub���Ư>d�A>��o�TQ�W,ց��?d+��m��L����>�R:��Y���c4S�7�31e��	V����fJ>�*�q$S��M 9
!�A1� ��ғNA<���CJ��Od�h���k�r��Zzj�
j�`��DB}F����=��q�6	�P�W%j	��?%Cr��⛾m���Pt�n?�UQ�Q��y�![,��aR��R�hR�E'S��9>gmD�wg���i�`�2=\_z��VD\���j�'��474���� 2�=Ĩ����V�7�Y����@���MIm�.��@6(���%g=g.�.��3'1Ͽ;?&�d2��]���?��1����Q�듽b��<`�Oڕ6(�6s��͚ �5�?ET�a�6�G�0�Ə�'"[��vb����7����Uh��Я��Od�v��1����=���i*�_�'�,9	�Ix��Xg�[�(ba��$2JY��0��P]�Q��y�5���J�8)�b�U�'�beJ�1�s�n��퉺ޏ5���/�/�3m������U������["8Q���	>\��˜ҕ�>��h�U�oF���i�X��Q����S�΢`y��b���毙"[� -v/~չH.�5�mZN�����i�>�0{�-�"�>'��&�'���Ϧ�ؤ� ih(�Aҷ���IB*��1�:���ޑ��c��Q3�X�����7 6�6pr����%-�
]e.���u��jK��;UA6١��bt�.R\�p$��i5�ct�K%�;���ř���g�,+�ѷڍ[�#J�<��,���/��:�(@����WE-U.<�_�^����7��$S�o�:?"��W�q���WI�h�=ڟN�:��[,;�Bw�QQW���eᗕq�_ϐ��hw�B(l2"2�H�wV�D�ۢ�뽬˂�湛�!?{��< �-.�N��d���8�<R�BW���f=�f�?exfCS�A4��Eu:��f�����I �y�>W1>�[r���K�Wqp?��vmm�����������r�\��::s2L�����ބz�9,<����\��'��Wg@�,� ےQ�!"GE�>$ R6l�)�ԿEf
���KD�֭�S�������v�Y�]��<2 }3�m替�HBP'ƅ �d��S�G{�����WO_4��RR+DK)6m5�E�Y��(��|g� {�4(��Ȳ_�b|,���Ow� ଷ��.���L��L�䝱��0L�_P�$6w�]^��j�;�ٻ,��3ċ2"#��p>�+ɻ��f����vS�B��/���U�+2�%8W��<E�CO���'�F�.��&�0����籐|� ��L�;�=(��4?���/����]����������R���,�*�6f_��t+:�q�vd`�cݷ��c�Xw�Q��`��.�w�A'�.6�p1 �8�زO��"((,�iX%��o�CKT��)!1l𿙉��@}�:�С�QݗP����|T�RMVJ���[�������ɇ��aU�pԤ��fK1�~�\�Eq�#fcMĄ��:Bn��_�=�VIe�h����Ϗ���`M�+AiBC�����E��il��[����ɛ�kAt�R�EwL*�w���Fo�X@�hƍx������I���d���ċ�wt6�ѯ�eܾ^�ɜQi�Hc�{l��q�W�D�f�J�`
<�)�B�=k��G<[Fփ��R�jVd�G� ���H~��9We��e[��k7����Λ7%�e�^Ǭ-1�v����Z$���#	^��=�����H�-�,�T�d���<S�ǸY0x���ɧ���R��H¯� ���|��,ׅ�������YE}'I�;�v��'.�g�A���׉9|��b�Ĳ��v��9"F��B���`
5�Q�έ(_���n���+MX��;�Z�ľ�����U��0��A�>=Ҁ�H��W.����2>�����p�����.����4Ǣ��'o]�l�+���bAk��(;��+�1�?y�|��ꊑy"o���RϠ����҄�>���$|�NR�;ٲ~1��,l����SX[�Q s(�K�V��YR���-mU������a�2s��v��K�S�ԙ�PX��
���'��Y�P;>�	`��~X9WF��#{G.��8ۗ��D}�S�O�s�����y#Ԇ�)9�_#B����[+��S�|�9;R��g8:���R)D�P��A�*iT!b!Zq��@м͋�y3ñ���3zĺ���w}	��`���no�"����%��X܄�:R]C8���7�:��`r���)M�\W=�W�nE<������U�,�Z���u��ak3�\X���;V��(s���9����Äw�t�����Q�[Gc߄ Q=z�"�8������7�ۄԄ������E��m���m�4�����N}Tkc-a���_�PFj`)^��.��-�qv�yF�f�/b�:�PJ�0_�qk醿�����Ŗ�����]�;
.��z����{l�,aL�O���
�� �W�US�d:���z�P�G��}Mʠa��3�2�ғ��mO[g�n�9L�4p�^���f^�K�����ܵA��
��e���T�nR�������<ZO��1�_�Tr���z}�L�� =i��Ns�������
���onPR��ND-��G�g���h�Eq
�nY��%ub�J��8�k����?UK��H'��Tb��
X8QR3�cj����(��'A�g��g�68ܯ�4
/��Rj�^���M�ܳӼt��s�I�/�/f���;^f��^������\-�N�t��\���`́�5�o-����pO�x�^�j��&��CB������b�����]4z���i+P�f�����<wXR�Ra-���	��'��wjfy?0ƣ�ݳ)99DL�KHbT��8�����rb�M�����M�u���LJU�u����j۶�;}6v"��]�zfzz�Z�Sn�q��tC�,D�w��	��\'�r����g=�MB?\z[����$c�#I�e���u�2��G~������ȅ���؊�eR]�+����!*Ϗ0TJ�N���O;�� �U|�!NO/V�KM�ֳ�T��?��=GԻwҨQ�Yxdy0�\#va��P�aK�ͽr����4�i��Oy{:�4��?�%�O<�K��:���<�
е�`�C'�=N����9��*(�����E���l���p��,P�oţ��,7�ι�~�>b�����%�*w����1�-�_Zl�w2�6{(_4 �u]J�.)���z֠l��#a��.����1%�	��Ws��@�R�.Y�&��?���&(ٓ�L3'���(r��r�c+4<B�n�����U�s��%K�:%�RӬ�Bm{�-�1
3�K�e���M�o�a|�Ɜ���)䜢�=ˌz��5ǡrv�ۦ9�v�7�ѕ��=Q��i�tIM�h�Op)Z�<�X���%Z��"+���&?J��<0�o���) ��:�YC�7ġ{�N_��Z������d�$K Ner�V�]���q�O�!���̒AJ.0Fܘ�Bh.ٜ�2_?s�(Z��%}��L/<�F -��ڞK�}6c��U6ѐ]�(�,���.9O�dF�Eޑ
��Rk�W^T|0��:��h�7��DK�Y֛y&A�V�D����S[��a(
G9Y�Z��cz����U$փ1œ�g��+���R�(�^.W'ي�I�׈�Q����&Ǚ�J`uM����V=fo��
�aN����'X��K��+��Z�4�(��]���W��2�z�5Ѻ�AŜ;��H%!0�C�H�:'����̂}3��Ǆ�ʥ�� s'?	�-��d�t6�@���ʕ�z�E�m|v�?J�]��k=�XE��gU����<�i�R�G	za��NA\�`V��}� ���
+B5�d�&�u��]Ϧ��Kqn��	�YatἤE񩓘�Ș��)� pxWQ2g7E�6I�_�?��YK��^)��_�v�N5�P���k�*�k[@�Y�k+k+2���9��S�z���5f��⾥�V�bX��Q��1%�6��#�ni"U�*��� �����N~g����0��n�˺K�w9!��*w����q/�<�&���Q4#S���+��0�Z|@PJ��q�lW�/�� �F݅�TA's���E�?�����s���Aa3�P�)m�{���E��]?�]���N��C@6�=�����t�'�F�'3Ꮆ�&H(dBTP�
���l���������b���@y�8���wgY�i8T�J�6 z0��x�����r�B�^�W%G�v��3�!XvݵW��W�U�G-'�"�y��W}�7��Hg���]%��0�zP�Ot�u�j�h(�S��� F��5r|�*���L�U]^N�:�a��q򨭧}M;Yw(*B{c���OW��l"�ay�+��W]zd���z(c$�|�#W;��3�!O��0j�ʏ��Q2���{�W��H�j�<א������1;J�jo�.�{.�YB���&��h�0e��-a�2� ��v=�^U��}��x#H<�V�Իq�R�T� �6�ul8��7��A%z2L�d���n=����-����|3۬%�M�x��:D�����8Y�(U�t�0в�ɑ��W2;�������f�
l�Z�(�����Xg�r��Wٛu1�T���|%�2@QdR����]]7?�q�N`SM~�-��wp��1�@}ݨ��7�����ҙ7�'��ב����G3#F�M{��=3��:OG�� ���#�>?��C>c}��9:���<k��L�Σ���|�B�i�S,�{<�G�_xMh9֍��9J�^T[����ɢ �`�xl�U�m�e�>_��MQ���@�Y��Z���m�V���f)EwE{gT��	(��n	�J�5�8&�~<����"�?,���.���'��ʦ	�Ls�g(�FqOure>O��{d�>v���އ��QX�5H$��'/ep���aη�b�%b.>S�.��؅�6��$X��T���G,�A4'��L-Uv�EukQ�Q��'�z`i�7t>� @����\nx+&O*�����^03ur_jV,�"1��I Oq�VY�L���B�rO���hwB����NLωsq�R�S�����s@.Z;\�C�ɘ�ù���-�$�A
���R!���dj�O@N�bIݚ�f��>�bsdJC����{N�{k�T��Z���cD(�}ޘ�;�����җ��a+&���b<����W��U��'7J6�Y�G����k��啁Wr6����,Ċ�DN��.�ߛg�Ӏ��=ߌ���N"-D�[{Ma�C8%�֟a��}�ԅ� ��-1^G$ɣ7u��@f����o'9�:�9iM�:}jk����0�D����!�5�7�w��e�J6�If����'�%Tr�2��p,nzzID��.C.��b�c�ׂ+%R�u��`��z��Ek����*�[�Q��!�)�yV#L(2x�	I��� !8V��y}/�	�p%\��W�ònT�8��$nֵ�V��v 76��Fʪ�W��F�?h�V��^/;�� �jܦ�z�����{O��Xj22�$I�����ZoH������B����o����.N��ÙD�,�w@�N���޿���f"8��OǾ@�Y|֠�^�}�4���w�����뺥��/f����@���Ev�s�!s����9�>����i0�a����5X}� I�H�a%��#A��c	n�N�C�|�P������}�b�?�G?�����1������Ɓ^����às����|���O�6tY@�#�FV9HI����i_
Pesed`Wc��]�JDpZ'��#Y
JqK(x�AYDC%�{�����υP��E�_�e#/���޳3,�����P_��Ҳ?Cc����`p��~�K)!�����zYF�YO�Ԥ��8K~p&֎�l�L@�d�K�(��s�"hy�?�F��P��C/�n��v�N�����������_`2o$ԯ걕�3�3 b7�8�?[���3� �?z�j�nW���g臙��ˬ^G�`�|�؄�E�+����Z-���I��[�������D*g���()�#�O�&�݂)LPV���x�����g���P��qVP��d#c���I�W1��N*ɔ�#������7��y�I��%q��@A�eɁ�8B�G�b3<���Z�N �����ot{5f4����d ⨋} (C��o�oYܜ��#/�F�VJ���&���W����K1�ﵙ@����5�8?�_�Q��0_+���]اc&���9�,�8�!�	L�(�� ��K�i��=[����z�8���R����X���%��7��3�V��&%8���I��;�R��d�şO�po�ݵ��|���YhF�v>�М �8��K夋������s,�K�����z�q�cq*1JKC%ߐLg�~���6�p�Ϩ��R�@�����m��K������v���եj8;�B+��@�aΙ�x�9pi��EHo�%|F$�Gp�I��*8_ſ�o��R��l��c�=�3*u��*�·��c=vY����^Ì����>�� #!+T��q���i�Ѭ�yvꤗ-��ؠ�=�W��T���#���R���� ��=�6�kB����9.��k��Y�v�M�Y�f�.�����_�f��F����9��x��<�:����a\����:�g��a,�9��ի�FhG�/U�i}K�� @`o*)D7�1����=4!�.!�Ҍ��_{:D����������V>c��	Y���/��������)gs�جPp�UI���՚5�!�pr:�V�_�O_��3����/a�w�e���T�|��۵�j�`��#�u���ӭ���>r�*�o���4�e��rȱ��C�h�ڈ������G�Y�����}Mz@,
NnZ�^D������,#9+��B�۱bi�RU����(��-���ؖ��<C���W��	��DG�9�ұ#q���}�	3�=�ش�!5Ȑ[϶Y�S����]L�o�y���y�9�SԚ�S�oQ7�E�'�%�M�p@��n�5a'�9y`�(<��pk"�E�<)�_0f$ښ�K(p���p�O�KE�j\Q�Lt�[n=e���&��\���J�[ N��4�%��Ԕ�S�����t8�U����+O>�qv���fXe����bȣ����K���D���y��*��Ecw�J�I{�yS���1g�q���~���fS�_)��q=G�g���3NPJ���'�9��tT�@2&���n�����Un���%��I�i���X�vs�jh���;�O%pG�+Nf݋�p�걘ϼ�#�����-#ò�H��� .�� O׬9���Ta��>������R�ϝ�����/�e�[yі�0����F���j���#(׆�
M�,��z�I��;晩�u5鬌�U䄮�<O�%s��AU�6�!)��5/y 9��z[{X7뾔���`nI�&��������e�<o����֍��8>���_�V�xHP�[�@R�4F66�A�ӍB:�;�&���h��-l#�H�¢GN�8A6>� ���rD#��,�jNT���I���N4%�^|���e��A�z��8���I\A��Cv��>D�+1�Õ�;��A�W]��TR���K��6�0�?��бD��=xe�l��m]��օB�P��/KP��~�
'�Ag:T�w1�b�%0_g'>H3�2���%�O�1���K&�`/� m���[��Y#�\�+g�B����c	O��=��c�V���	�^Q��Y>��b�opOA�5B�6w�����p!h��/EG�i����=jeDS?G�������ޭcŝ���wyw�Ȯ���di���@HK���69�H�߰`�<uIT�־O%p�1t�LSys�NM��n&���>Mn\,��Iw*"\E�}����W���Fy�=4�ώ�� ��}�\B�ެg�3�UNZ���������s�)GtL���&��� �'��t��*���Y9�J�R��.�tI�Ԙ�W�WGF;���(�Ն�(��{]��z́i�y@O�hd���}���z>��u�9�e��%\T��Q�`���Q�!p`�Y��x`��*�B�t*��qó�D��wh��~�|q�5�S��ȿ�В�M���#��SO����i/;�H���ec��d�V�|�A'�k��IL\�$���k83���ߩ�p+�;i�`ا{7n�1]%=t4�Cc8B��M6o#?ڿ��:��PS`/DY]��(z���s�bWz��/��52����6>�Gx�"��l�`A�>)����OA����L���5�RI�=��ּ{~�Q�R�C���r�"��S�%ډ��k��Hh� �R�?��b��r1� .��#�p���؝U�����(���?������`wz���_���&��a+i3���*4�^���O��5>e���>c�.�,�&\w}�Mm�xn�k�#��3/����W��sY��UߪH���hj!�����$5�R�`il�!HR�HhX��Y��hΟ�~O�����I1�F��pF���)K�Z�4�.ƥ%m"�*�*������}��P��_��@`F!�[h���V�_��m4�} +�2H����P� ����^e�?	3��K��m�2���T������$��D/i�6��'0��B��a�fz�EDʈ8���e"7��\�g�j�W�TV:6Pe�#�/�B-���lC*��t���<�r�'T�����`Dۯ�A��A9ۻWx?5��3\~�>֤qn��F��r���g1��ϳK������� jj��6ìߺ�t͏�Ÿ��[�����O�{�QuH��d|�b?؎
��%��̦�Mm6<z"�RDS�e�i�&Yɕ�{mU$�u�8��ΌZ4��U���	�t$[|�Mr����tx�K����-��ު��DJA��50Jmm�-��?i%0w����ja	l)1��ǏG�� Q��O��b�D�l;z)�A2Grs�p6E
Rהℜ�|�j�k(��M�D�����S�Ü��-Q�ۉP�%��(Bw�����c ^f7��6��yNt]�-��_��w��WT��p�hv�3�֮Z|��$�����_v�`�}��p���=�;���ēU|������	<����F����(2���������w&�Jr^����V۾�0���-��G4!]�-K\xt���������T3��N���PL��NF�R��w,5r��4�+�-�Q�"j�68%�c�ɮ�����h��J8vZ��$���	f�;�՚^Dt��G���<��2ɔ�h�bh�wX,A��S�aFC�<{�9f�̞��Q'�`5BSY?�hf�Z��z��Y���=-��������Wف�H�@�����wIB���1ɃAS�V>!�st°]`� �\�g@���	�_�HM�BY cKS �"f;�Y��膣����+ +����$_�'�3���\\{�� [jW���wO�s�����(�D�C�x��Z���i��YL��To/4b���Fv_��z��s�^�ϒۮ�lX[.l���tO������0~p��Öy{�}�T��.]�=	�?�=j�U�I��l�Z�����B__�5S׼]����l�m:�,e|w����+�d/�G��K��(�W'1�bH��K��R���[F���hc4O0j����+�a���)�z��(q�U��5��v
pb�_�D�/��*�9�7�YVU�����o�r�~��5�r*J�� 
�����������@-����ZP��8�sF�]�@yFrDal���a8��9�ʓ�A3�чτ���εC�%�V�=[2䴄�_~Iш�T��$���$�4��B&]�/Љ?Oh�_4����JO��7�)-�%i'��F���`~�������~�y�o>}ɫB+�aJ���Z݇��-A0Ϥ�.���ĸ ���</�j}	�~Ƈ����'O3t�ą���|.���	���&� ���6�����n >v�U��,�����{��E�U��6+$ZM2P��L����&ިi&�lRiS���σ�F;�4Ř��[������-0�"�mH�'zˮ
̭&l���|��-�a{��|�╕�0��("qp�dQt��*zT��MݑQ�H�H~��&��#�z~>ӪSP9q[E(�S��{�>i�4�Y�X���l�"c�c�8�+}(�o�iK����T�Pe�R���lV�[ 0�F�gWAE�T��,�5��k*�]Q�=1G���ˀ���S@�dF�7�~�S�(��<�`W�g5m���J�^w�(s١~b���
�n#��ӎ����:���ϭV�H�Q������Ϡ�,m3��_��D�7൧xV�պW��Y�	P?G�C���˭�?Yh�s��{�0�(���:���o���J�j"��+`Iy�U�oF�_(�rn�#���>�����Se#�L1?`��kN�0q$A(��#
��GR.����D�-���F/-� ���%-��^�MTw��=��H���>���ƾ�&��^�寨�+�/�usV�M�,c� �D���Y�"�Š��F��9�q�r�ϑ̈́3%�@�s�/��~��ޞ)Ȣq�q�o����^����$fI���܋	�%X>%4� 9�v�izk�K�(�}j��9:�|���}D�����/k�i�����fo�!��uA�h���;���e`�7� �㍻:���+�D���P=�o.�׎n�Hy���W�ǰ�>j��=Q6���4xs[,i�Ԁ�؟�����1l!,��wV���Cɚf��NN��R�C@���n+Y�|�ؖe/Ϡ~��\c�q�3�A(6٠��I5�n�p�fU�%������#�&�Z\ȫ����Z�WU�.q�����X��;�#�E����8��En�^`�d6H�o�pl@��ׄ�mLP�t��ƥ0�;��U�����ҽ̇l&�8�+48[��|�"3�[m���O��f���H'@f�"�EC���c��I
,%o��m� �О{�ȴ�2m���}���|�p�FUr�!.�T׃&W�P{�A���1pw;�.���cl�?�r �r���UG�zO��.Fo�s��uQ :���U�mg�i(�g�I���', ���Gn=�4/��c�_�O�խR�2�5���ze�H��v�0��3��Ҥ�Em>� #���r�A2��تI�=�m������΃�s���m�l�(UԺ?��r��q���_'�n$�@Lb�=�i��@�P�c�͖1oI�%�3��l�uH�R0�Ҏ���1��u��{9���"�T���w�sy�ԖB�|��C��F�DL#2���A�
�{�cD��˶_7�J��J�LZ��կ�t�]�E���8'k���� ,�ۑ��p�ϠJc�v�f�g:��f�˺^"\_���P	 �x�#[��k3<S�W=���`�U�:yF�a=|��B$�:�}�o{g{�2_��b�3��kؕ܄�x�N���f����A8h��gu�t�G�
+i�|H�����Y�^�9G۠�{I�����2�YX<Kv����G_&ZII��&�l:�UZB- z
����Ut6��Ro��O�����v�G�	��U�� ���u��t:�(��į�Q6��C�����}����Mg�dԆ�>H�@T-i���7���O[�>N�J�N�9ȾP��i:No�m�����:��`2����y���cv�2wd����aH?�"G�nUG�yp51��Ã�wQ�%�m��,��:�a&Z���:����&V���Fn#��8�t��S��I��)�4�672�??
���҇b�K��r��D͉!e�t��k��Ct��[j��\�Y�ƟS��X�d�Q;�!��c!'q���Z*���3r^�p��4a�C�������O��W[/������*��m���qړH{GG?qDoh���F'��A1�P:�B�4��ꅌ����h���Ϋ=�y��]���XX��(�߷V�b��E��g���=I�<�g���F��� S'��>a�^�I�j�$%�b�X��5�����"dI�I�{��4m���'d9��	P������,�t�:;[�V�x24��ڑ$H�Mb�/;�O͔��I$;^��l��{�� T,��4v��@�:3�H �j`PD=�i�d�`D�F�C�'�A�c�Q�]�O�=��	&�7����c��#��/'�*��5z��a:����=�7�����=:�q��
��"!
����u름�9g�c{�31S�H�l�1s����r�oF�����2�n�c�+�*��X��s/�Ot�����Vt�噻�҇��� ?���spL�=��{yizl8i5���|
$�a�C�}���h��i�i�u�1����ql�Cǧ�����Y%s�����-?�ڈ������ ���6�pXkXƝR���Ρϑ��6��@3a�3U̐���ە�m�-��ӝo�Ȏ]Y/1���"�ʒ��]�o���8T�����
��B
����3��9�-�Z\�
&�����Y}��#܊���p�/0�p�2�
��NLGoD�bMe�Xi��������(9J�������bu���S�~!��*����e�u=��HV��`ip�����8A�}��[q���Ѝ�
��A�<������ZGr����W�؞�;6ny�_�feb��M��"�螆J�A΂�E�F����o��_�̕�P�}#�>� �U|�ZE��)�)1�#@Rv��v�Q��6�˴A�ޅ�����و/��ȁ��K P�7�7Vr���Y��%�{0H��̋d��lJ���1�Y�c��۷��د}���P�A�$�<��=��V�&늛jaz�*�IC�hj�-7�<AM�
d%J����`ax�eN����i0���$�!���r��f卍r�d��tR�W�ݵ��c�ndE ��skąo��b>���
�;��\�L�s�L��9]	w�	�Ou��-א�)�Z�p�?�V7,�2IZ���ĳ�vJ������/M�d��n�n�T@6��w|�������f�F�t���z m!欸'�-�������u�;���~ץo�P5>�3l'�&I�V����Z��^� �ёy?حѰ��z8�n�/\���p���`�o��7 *���R&X�ړg�:�_��=*��ZI���U"�xߥGoq{G�C1ǅ�wX����4������F::��=�ơ��s��o'���h�����Z~�T�yΈ}�=�~��"����m�!������&�o4��и˅��7��,¶"`pj=�z7�&mv�Y���/ˬO��b��n��>��O�[e�l  E]���!`*�i,������xĚTc����Ѵ���o����9r��'�֞7���cL�VN��X80ǧ�g欵�k}����	��LO���:H��gX��%!$���� L]����H_#�\R��)l�N���񉅶�cIv�E`�T��:�(�C���"�����4�^�H";��ap�����M�p�6�](��~^�#8j$ˠn̤����­|S�����D3���Y����}�{Y�_X�`ꐋ��M��M���=ЉJЮ?�;p�w��w*���9� ���e��5��F�*��ҋ��|��݄�W��ݑ�b�佫u���Zɥ��gP���i{'	�����q͇(.HBNO���}ۀ�C�}�]W����S���m �	K�x����O�a��+Y��2.��:�b�0n� iXJ�ȁ�u��h$y��Iq*o�{�o^�;�p�Է5�o����$��R_��1��g�!l�j�G��I|?�V�3ù��7( ���gn~���rzr&̸�cռ�k�̛����0�y\]7��ή#*�}�lnԳ�L�d�����~W:�(�7g|[8���֋4�ֈ&�q2a��%�񂢁����/���%���ME�.�='������j��~�z����p���	^���]�r8��DK�����o~ ���e�\�Ĺ�� ��4�T,��¬�޻;�?j��?r%�!c�Ć�� G�͉?/���r�0=�������1N�����Ħn������'�*p�t�����k��1���8'Ӑ��vف��[%-��g��6�Lm+j�B�C��˕y�n�b�ۃbc0~2G���M��ʎ�º7/KW�H�5�����;�����&>��)- S^ݘx5߸zn�uB�G���?�j��J��ۊC�8qfU�p�~��P!�����>�E�$�,Cj���l���8ǔa]�,����:�ɨ��AEE��~��'�lĥB1f[3��3rd�ʇ�@��:"�����d6J�Ω��?]���D�r���O���j���X}1�<n'���cB�d���{�^�_�k�u��� wKAV�{��ׂ���f�0<�ߠ7�Uç��y�z�⠝�ڣ�3�v���ÿ�����:'&`���,R\Z��Enyw��#�v��;����=v�� �_H"�L��E�$�)��7�v���A����E���+��0s������6�{�Ajt(���`h�
�,�'�������H�8�U#�S��Vw��{/������Rpzl��H�p��-,���H�x��𔌦y�G�Q&�v�0��t���3]�	ho�Nød��N
F��nit8pU�J4��j��`}�F�{d�o�y����M������/$^/��.����'�͝y��ٸ�uc�u3wvV���3��W5���(Y!���"��7�N����Ņo8
bk ^����R���V����Q�OOJ<�_��&0?̺����λr�|�82��x�h���'<��#��s#���M܇���@(Z�|���!y�6��ְ���^r�{�2�0�,�K�ap�3iTΝ�����:x�D�t�����Xlz�RX2^��+1�?Lr��#ܨ=:"�0*"R��O��ux�u�J+�µrg%�MU�����T(d��d���)ps���|�e�Qߒ�}��}���x�N~�Tq�x%#���*����	��!�x��̂������fس4Ԋ b#8v���=$Q��͎�VŨ��ً��e����6��)@ӐL���"����'�~��+���r	7��?7f�kGڤ��4hw1Ά`�����,�y��`�;0�!����;m��s6q�K0��0�L���C׺DxN�C�0\J�m��8)�J�����s�"��$8h�	1e��=���1X�m��������;�ӟ�߃+o�����Ʀ]]�Y,[q����n�x8t]�b�B�����^XD.c�_.D��2��gD�'hk�_���(��~A���M��	Ey��ܺ��Q�a�ɫ� �8�� �{�{�ݔ;Y#��[Y!5 kԵh(�6���(�Lk�K԰��\2'�ƒ�_�e�][��=X�K�m+�;q�
�o)�QL[,�f(����ƽK�/�urLS(��:pGs��q�U�1ߖ�N��E`V"˯�7xܥ���({��ш�C���Xl��-\���)3\��-���sѡͩ{T��ŏ���.�/���額|Ts�{yh�<��[0kDk� ")Sw{H�I���7bb�O�y�d�gҊ8��T��]_<)?�|@��S%@�O�f-�W[�(��i�����[��b�6�~?��gJ���rKJ��¬ �|�v�7��V	�g�ܷAJ|�����������`�^e�$e�$vA��SyY�gd=�{}���.8g�5�pN�T��Ŝ(�"�e-8#X�o;]� d����ȳ͗�������y���D:�:�n�8�3%��x����Ӈ��Y3˒�̀,�SO'���)��c}������a�x���p�*��C���~�.&6'����'W(��!��it�'G)rp}e(s*d�{j^P��=�������@��PC��G'�b��N~�����H.J�֣$V������B�6�Y¶&&�p��$�H�l�`�A��<^��` ��F�����eΰ�d���t��~��{�-����*kn�Q���Yl�`:GJ� �1�lje���/����&0���&ު��Z�.E�h�w*�s�L�u�:PG+K��qm���]�n��@�`�|4�t������jx��)m�qq�p�n�;�e�ߥ%��rB�����Hw�ޒ��O���?�����J�ݿ�U���B�<�r�O|]���&b5��TF��)WrZ��հ��b$b��������̣�Ni�ɷQo9w�k�I7���A̶7J�uLW�v$f?��6��k�QF��o�8��B���U��Jxb�Әk�_����d��be!���_�!q�}FS. PNC�T�Rqp���(Z�b��H_
��y�O�_�29��QU�wzUB��֠�VLJU̟�Μ.U�d��f��52@��|�BPS��l3a,=aٜvؠ\F���H�-�jU���7@�Ü!�"��5��Y��Л�Om�߲�l�un2�T�m�-��|��H�����H���D�%��}� M�i�0�h����(Nvu�H���sp�R[�h�����Sߡ}����-�鶜6ߋ@���2�> ΐ�5��k���z����Q6��UCm�]�3���N�@#�sa�����r5��N�v0��nPV�n�\���ӻ�u�	E_�"�����i�HJ:e�~�5��ڼ��qE��_`��8�ק���q�IJ�ɿ��=bv �I=%���)D�K�N�n+��R�EFJ`������L��Р�ٜ'�[Y� �u����Iu�ގ�##-.�L�g�D>���	�O|�ަk�faK*���>��:��$8��|�Ԍ��t�!����Ad��;��'�9K�?؄I~���
7�!���9V�8�����U���3c�|��8���і.�2^&�q�,��ޭa#Ln6��@ n�'YW�����!�M)�'������H�y�B�5��kv�9Z��,ݴ���昿�E��3�-��So�0�c�(D��bi�K���u'tg�X�@�I�QqwX�;�0���B.�\�a2�"�� �C`S)J���ߪ���(��Q? �J���u�.*sbpwA!�0�!lNh Y �
�w�8% ������݄�Rnsx��t{'�~��Bb��9d][y���֯Ah��@9�G=:���<����Bf�Y�	-�5:8�Z�vd
�E���)vC�>���a�]�u�������!}����!��=��"�m&��u��g9.d�A�:LDAv�H����"�/��h
��H�}�i'���{2�#YT�Ԙ�;d��{�h��05������#���a�,�Ut��úk6dṐLLaey]�|)���Pt��ƃ��1J�)�G}\���ܵ�UH>����
n���U���$�G�f�k�0[��OmH���t\q�[�Q[tT�>��j��U�}v�m�lL��CnfqF�s��aq��~Et���,�2�Z#�1_x����C���uz���Κ���$�g��X�����J��w����B�����Y�-W�c^��JL~������~YҢ ,�� E�N��v���|e���GayXֹd��G_��d'�X8=�.��C��? �=��`��f������{��IW`,���K��~����vۗ�x:��c�+?�f?F���c;� �-�2�,�"�yU+q�3�L�l���'.��x����ճ���Nw� �î�#��rE(��J&(�hx�c?,!�2H����.�f\��"�F��#w%Y�ת��P���@�U�$I��پ���/B�:���x���m�K��a���$�Dr����]�� �{�3{�\De�����`+�䗤�ʘu���x\��*IH}��l�>���2��&&�L���[*��\���"ӏ��-�p�6j��s���I͖1~ q�t��Nd6� �������}3���&ՁBU�jE@+0)o���6�-�;�^G�O]A�$B?}�� ��;��f�v�o��y
�s�}9z[
�X�g,����V��VV���c/�y�CC�[�@�k���/`D�#��xǱ����/�:f�
�,�9������C��G}��6rY���
7M�
���[irO���cư}ܻ�Ae�Ӷ7m{�C�0����Q9�l
�$�cDSH����Őx���\)��K����{3iH��S��ˑ�S5ff����,�)|�n֮�[n�~@[99(�X�Pz�ǈ��{{Z6 �eo��F܇��j��^��><,���J�-]t��0;n/�һX������O�}�6{;�U�.�~R�Q��)jyx�o�O	�uzO%�����rj�%���� Ye����4K����7�C�>�C$�k���ޒ*gջt�LC7`:���H]�wW#�����	�6���U���Ⱥ�n���!LBͿ�[�2��ny��h��@���;M�(�)`��:�'-=Ez�U��EP5���_����ea�p,��B���2�S��E��L 1�����+�����~3B}�HOU�Z=�R�p4Yv����6�`_���l�x��������b�9��'�v�����[N��SpT��_�)0����o�λ��P	� !�3p�YSa��;~�9�n������r�D�?��r��|�7Ϋ�o ��L��&m39��TpM���+/�x�ӡ���|�k} ߪ�9*��6ptv��-È����f� ��M5&��zu�G=�o����ݰçD���[w�7r\��PV6�T��6��0�S�]����E_ˣK�_$�x�)���B4��~��[w�S�`\F�_��b�vm �Ui8���d�t�x��ū��g�o�
��oWF��$:h���׀��[��Kuay�a�AsPRX���y�"��Ө)�*4��(��]q`�B�(��\놖x*�j皡$�Ƅ��l�t����1s�2�%@e��=n���2vT��5�J	������W�`�����  ��=幌4j��P�����B��z7��j&z>ճ�53X�Y��fU ��~ס;>%�A���k,W��[���J��|��;�puǍ;hd<}�?IT��$��E ���DԑΒD	��w�ש�W�<�Qsȕ��] ���sA�d��_��	e�n�Ot����n���ϼ[?!�
���s�j�ũhq/蓯e`:����<�3�v���]�;}�e�>��A+ŷu�#uca
�/�K�Eɑ�)6�v_64�`H2�����j�i��'d�h�lwWwa � �%�l�99�$���U깪�	�f�r	괧$:31��f����|�3*/&�n�p��+di�>�*�Ƅ��O��ś�\�{�+��i�;�3�#@���~�j����%��'��v!Ož%�Zv��3RL��]��-z-)-�-�Hjx��l��ᛉ�-;�\�Cucn�7�҃�8 �v�ӎ�n�Ɩ1�Z�z�z�Z��6c��*�$���*n�?p�?8��\)6�-A�:V��-�����|��q��۞PՔ�;/�Gei����ۂ�G��د�ݛQ�!C����3�%���ߋ������bp��*�f��I�0_���/	�ڋ"��
��r�BXd�����Yo��P�JeFo�.մ�I���j�`qS,�4�Z�t��_�І���q�,wlM��Ƽ�Fx��*.�Y�u ��(��Wb�a𛴨Ƌ�v�n^(끖Q��x�c�B
�СMΟBRY_�!{7�Y1��%d�t�tTp��SA�?�`���&��.E|����A������Y�����3�V"�C7��jg�������k懳Sd��!��k'xtbX%��Z�񉯓"Eb>�O9bH_�-�X��s�Ո�S\F�Հzf#�@��%|0��\���[E9�x��㔍��o��5�ֲno��~܊Mq0��%����"�!}�!?aV�\1�!y�s}��o�!t�{���t�z�l?��3�3� ��T�Ȩ�b�7�D��e��F�mźֲW�"�gWɏO$��u������8h�}j�Y� �$��"�ֶ�����D߅u�_-�ӊ�EV��@/*D͛�i���$�;:�Qr[�%�#F�8;5�����2���-fB�1̠Q�*}����'�Mj6ЅR�c�R�\�����7LX�F5"p��(�9��Q5F��J�r]��ǻ'��!X�vnX��x��I�r����G�<k��G �]�"AX�����m��LJT�a��q�Kߨ5\��^����:�w
X����(84������D�<�~�}�&SQ�V3@�x��%pޅ��?�&�������*�gƐ:Vw�g
!\����7U~�:�E��A���ܙ�$ɢh��n|�� �Δ�8/ �;�\��?�a�NB�3���1q_��zu��)����e����,��B��v�Y<������J�v��V>&"�ж]|��w�zOTMI�2��V���Y��ɛ���\G�I&�2h!N���,t����@�_�Tb��w�������G"���15��F��A�+��I\>A��_��X�s�mI���ˤ���e�	�O&�ɩ#��	� k#+��:�sn�,݂S��m۸��脼10�P��Xc�2{�Z � v��'H��L���p���� �1AXE��H�v=��l��r�S��H&F�;B3ʖ�w�#���I-݊����'^dZ1Lj_�C7?�X��Ɂ��4)|7���Ğ��,o��󑱆i����k16��*�UT�EItף�����}w@vU�!���AA�ձ��/���V�,�<:��]Ո��@��@��cˊ��O���U�Á%�X˿���U�)P!z"��� �$���&"N3bQ�:������$�r�-�/��
�F��L1���?y'�r��-b�`�Qޘ��AR}�a��+e[)�tO���� ހ��0�X�܋��>��&pn\��}�;u�ž���D��ڡ`{���C�U�V �x�M"!z�&��{��p�}0Q����G08&mJo�a*�!`�lb�8�ǆW=��ȁRU|ԼG%hc.	�.:ੜ�;�MƄ��/�A��^Z�h���N�+�c�k�����K%��U�qO�P��B����E����e�,\*��$���^�M���e�2;��6�B��@7�b�u�+4����h�P7��bf��Jש*�~7����Ϝc���F}�ʳ�%;U�O��z��*Es� �4N�����+�n|g�C��|�Ǘ�W�I)h��YM�kH1�uX���J+)��sT�ZNx��~]vy���h�H[�ʝ@76���5�,�"��a�B��T\p��m|���eo����(����� ��Lm�c�v�L��0�,h�z���� J�D1%<�f�c(��jڙ�Y"������!��W�� {�NL�{������`�H����j���A>��K�L���ʡ���R�gOG�/z�0߁�����G�N�{���lA
����P�7�d�o'0읻�s4�L�h@%���V��o�
/�U�J/��e����&���oi�(^���o���E��UF��&��h��E(���=�D�ڡW5�N�Fƫ`��hå�kJ9��'�W���eA޼8�r�)�6(����D��Vs~pq�Gؼ�b�,v��Q&��Q|����
���	¦�I�RZ�����&��Xn-�
�	}��ھLeڥ��DTm�Ϋ��d0�И<�oH>ۗ�w rm�j����8�88��9�����)�zj� K�W�Edհ/n�qPD��	�-���g���-N�Y��<0��(���B�c`��"�YR2���Up��U=n>�Z�$�����0��S�=����_�#�T�b�L�4FI$�p1��;�ΐHh��,�-R3@��ډ��rD���n/��̫�WzV�(r\�� �` �u�|���:��N��/�%J���A�-�e��I2��rG���qx`�Т�D<����i�ٸ��>�y�¢���s�{�g%c�gو�J��RA�ބc^���ωT�YzQٱj^�ͩ�t=yba~��F?�k5�%靈����l���O+B���1�}Ʒ���6�iP�����n��8!"���P`�R���SxJ��/����ci��q�^�A�+�RZ9d�)F�F�p��2����V�S�^�p����Y��`P��|D��{V�������$�Ub�P�w���ϟ1�8|��w������ι�SnHi�g���&I��i5��f��3���o������$SɃ dc8�A>�az�����yIKVGN�~��DyG> �FB��)�����Buroq>B�l�S�5G�����yٻmt\(�t�|0�{T17�Q���G��8�^��Z�}�d������ʈ,x���G��ǣ���?	�V?|6EA��S���R�rTr����tP�]�o�yǡ�K�)�4:�r�|s;I@ET��Ypb/-�1�*��ENڊ����Ɣ)Π��N�Շ��l�8/2��:��F��_��������o�.������§.[������*{�Q�^yӔB<�D��Uv� N�� 9v.�=��h.��jkX�[�8�ُ�V�c*���,n	��p�	��B;V�MNfl3Q؈bzT�`v5����!��E+���z�pZ�u#[˫�R�^U�����W�e�m�IW�5]���"6ٸڣogOI�f��9W�N�	���3kT�s9�ٗWȆ�R1��8��p4������AD��鍨��v�tL��y��7WIy&�9^�Tސ$Z���61�r ^�T*d�wA�b�I��.�3g���p�m��V�@�*t__�D�bN�t��>a�L�L@?㕦������ْ�j3\�b�r��fؐɳ6#��>vAϚ�������a�����y~מ+��*~+����BM~LF��ƅvZ̐`����Ŕ�@�h �q�9�>
f��P�]B {/��W�n�D�|3�Yj�:aRo�w�
Q��I��	k���s_U0�rݲ;;�XG֋�雷�j��x�ͽā�����y�����3�w���s���@v�cƬ��x����^W��c�Ik+�n]u)!������ѩ_%�-�g�bX�+�x�#A���T�2���2��<r��}����2D�)"9����k�i��K�b34	 �p�5W�|ǚ��ڳ�I�nd6�����!S��3�����b�"�OD��v���i��c5nRg켸lŔN:�ʘ}v8��:|��N+�@p�M̄D���h3\��Z��r=��M��k4��
Hr��m���%Z�%/����rJ��$��s�D�@�%�s^�z٠���-3�M�$0�k4��@sn����L�V��1�N�V���y��t`�)� �aT���2p��Lz/2H�Ϩ��'ϲh��w ss�k�W������G��?H��P���O��x�Fc�>����D�u4���J�flF��� ���D���f(�Z�D�%��Ȭ���nn�$�oSU!:<��+���6L�gtf�屳�����0�<��t�Q�C@�B$���Ѷc��P��:���E�z@��!jh�7�PS��$ù����l��"tc!b.�����k5d��a�gU���^	�~��qm���>��B1zz�0�2�jU�����?�A��V ����0�BApV=�0�YR���z� ���A��'[~.U��
l��c��k8.�(LKH�������f��5މ���3�/	9f��$�K�\�J�w|�N�=U��2.�}���qV|���yxL�Տ����@b,��vA�H��*!�����q�0ևn�R�g�X
�Ft|5@�ln{J�q�.SK�H��y��}n��Y3??�D�l����i�wqN4D�lG�)���� җp<���g�F��N��{˥�^�_1��6i��M1_��mu�Y�Zt^"��n_Ղ���kǐ��f����H��s'=��g��S��P`R�-�l/:��f�ʍ�e3ϒ+�r���*��	@�C�Rl�i�Yz�Tl�(Ś��>����goy�r9��@v��Di 1{j#�<�X�ǘ@���ite�N��j`{C��~ǔ3�~����Q�� ��I/����<�4s�G$���ƚ9_CE���b&�;̶�0
�֍��G*���r�;�)a;r!\`�U0�.>�9��(�8i��ʠ	��"Q���7�^�x�G�����~I��q@kЎ�%g�#@�#�4�jު��;,2>dQl�Oy��z�E��,d릏�L-��yj�ϔd�P	2��E�S6&Aq�P��4Y�L�����dh������\Q�������;�z�e��@L��%��4���0�<�"�x�	Ο�i���Fc�*�Dk0�`��(�
�	O,]����3�:m->�l�Xل��mG/�D!z�g1b�"��+���7W�i�g<�I�n ꮏy��i��7/�MN��v����]ު�&0t��6�����D�&��lʄ���u�;f�!$?(�G�@�6�pM�q[�����E*�N����"*��v��[���h�S�.����6�LsYi��s�q>5=��hx�e^�Arux��Av��In+o�^�=}V����!e�$�T���6)��"��?vկAN&q�'u��a�չ��%#��ۻ�2��)���m�| t�9j�e�A�]�"#Zs!�+��P�s��d�[��yqw,�Z-A�zR�~�ɬ4�J �x3IV31*�00J�����4$��m��a� -X��y4b���f����0Z{�:���x�"����\Q;M.��wSh�;/71KP���n��c�z^$VT���H]�3���k���X����ɑ�Zg�~N�<�����mEq����.理V��І���
��t=�C�c��x��V�h�MY�����,��L�q�=@;#��M�50���l���n�k��F"�F=��Nd�D��ea�NN�Sˇ'���)��/�a�[P��e���-G�(�������Y �w9#��$g
�%Ʊ6$�GF�w��l�J$|�a/Uo_�͓,�������O�^���*f,K�"y9�\6���v�_��c�y��0�7V�����J�rQ��J�/��l�� ���B�_��B��>M� م*�M�o���7�0uW�1V��K����cWg�[)f��T�x��^�؈��RB' �"��u.����� ������}\�~��9�9��;���`2�75����r[����>�s{d��S���Ɖ	`�8�?3�lr#�S�R�x!]�ܐ�S�kҢ|`H�vab�`�F�[��3Rmm���?��6��;���v<r4ec�i����Cg�Y���59�x��VA}VW��^i�&&z�E$ E���������L74���a:�����K�=�t����ʆ�7*��z�Ǖ���"��Pe�_�e���	i����[V��^r�mNn�3e~��j5���K��=qW��Zm�^�w�- =�^��&��>k�Sd����g�*���|�i�$����U�,��b�䁝�1~���9k��2^��!-}��i��,�B�l��y�by'iPp��Ժ��z���+�۱��	8�{���T�oZ��aea��~����'}�E�	E�����Е�ˏ�jL	��Ǽ��}��)?�����yR����&S������yXY#}�R��b���G����,�LS���T8�_v/2�Q�kE�-���ͨ�r�^`:�w�v��R��?gRp��"�ޯn��T0���V��+�V���̒7��Hv�p��?�*k�S�y�;o��<֒��3A��Ov(���ҧ���o�.���)b��T��bA��x����	=l�����ږ)/��W��/I�(sUo���eU6�����/Z���!f�� d�lh�x�����D�������O��lݺ!�t�3]T�1�= ,]a [��h�be��'vؑ��ڌ�}��:ݺ{��N>[ �S���ϝ��}��l�	�ܮ
����u_�w'�<ډ,����f�TGv��Ӳ���'��&<�]:<�Z|��"\��}1�v��N6ϝ"Ąr���ת-^�`Bď(Au���T��x�h8.��~bݗ͉�9.�Ȉ9 ~������!�
7T���
��6��e�W�-}�H�9i��n��_�������3��C��/y�g����a+3	sd�j��G��*��7�ۡK�$��a|��|���)ma��&i��-M�:G�#�U5�-A4{#�����w-ܭq�8��hU[������ysXLӈB�{L7Do.���,�����fq&N������z�]�-��B�� s �ǲЍhH%*b'�Q^.	-�L0ؗ�d�+�@��m�:u[��3���Ҥ�K������'��A3L5�l�5� (�VnGö�I��+��6��.��B:����e��1!V�%\!^E�����C�1��?%�=6�"N'e] �i�L�{������`S/�k�{Q7�J:�\ wgQU�!��y���T�̦�"�"���C��x!BSQ�!�:��~�**��\��[�qI4z�ߑ�om�����m D���A�C�+m����.o��1����,�%���w���귩d��C�z�/Ė��^�]z�|3a����d4�i�t��d���=H�3��&	��d���f�B���%��|�>{���O��m�[9����V� ��8Gr�{��d��d
E���gQ�T6<ŽH�h&נ1�։�qQl�W��=&���yZ��5f\���iC��H�X­I�c�؂$:���;���Q���|��{�h��9�����O/���# =RR\ ���<3�Ǌv�-#h!�Cl�<��a�߂pc{x}gzu�.���Ĉ^�]�O�_^�
��_�-��ɬ��}y`���8���=��P�Z�1\������	V-��|O-�DfF�6�m�B�K$��������;&�
�X��C�{f�5�R����׉ڕ5i:g�d����GT�"��9gi#����%ΥF���>%h��i[������/P��܌�\9�|�kf�'���&��W����h���-~e�����W� ��sqv�i�>G�� PK��A1�s��JW]��\B.��i�����t3#T�ZG>���2߳>�[DΌ����]�f�1H�"�Se�hcP�Hυ�o�R�ъ1|�����0�O�u/6׋Fv&�����w�g���k
*�*Lg�U�l��Sߒu�M�4NAw�
b ,*č� �[D,�hB87�yO��m�1�����h�\�*+1�9<��|$:��X@��o����Ď��;����tt6vN��F�7~�����:���bɇ����:b᫲�UQ\���Q��
��N��9	cz;',�:�%v6�51�{Y%D~"��̋�;��J�ݨ��>/���Q�_r�ڮ��K�y��6(���������s��c�7��C�諷���3]��G��A����
��!0�!	S����8�'����S���}-H�T��q�k�y����Zw5��$��W�%��ͅ�}��l��� ��ڽ��
qw��X����a����}��Fbnp7��h�Ǚ�uq���:�Ƿ����۷'a3TF�����ޓ�&�j�0�Y�3�p̪���n��\����u=�aퟠ����@x��� �xLE[kH_�`f7.�р\E`q
)8�s���+E����9������'�L�����/��6T�ı�;��Ѫ��1�嶦U����n6X�����#\%ϷB��R�µ�.��k�nw5f��$}a�B�Ԫ&Ŝ��/̜�E^�C�ԷK�pk � b�N�߀D������_Ce�%^�`3���h1��dY��qC�5ܩ���sl�P�}�tr2�$E��ɉ��T\���@O���x�Ms�ʃrq����E��e/6�abD%����ƣY�X&UrY�s	�C��rdW���<U�^�)��D�	�_΅Р-�����DiQ	������g>�����5K���0'��z��~�/o�s�����ӵ*�8U~gyo���2�ɬ}�����e����wH%%��UH������g��o���܁TY����n �0�7H���Bd�"W��v�^a�����L��͉�2��DT�ޡ!Ի���T�[E�c�ʥ�`g�<�w5���5z�Ơ�����Í��C|�F[�����q�u��t|�l�~&�F���(�%N+�k���\��> B�_:F�+������-)�3Ĝ�d�������#��A�:��Q�u6�܀ӹ�����Y�ZA��k7��	��K�CZ�P�>n-'��|��;����ՊbSPۏ�w拋�;A�Ew��odk������C�5],��X;�_6�7N�r�N?��R�� <N|9�(�p+Lȶf0L^���MQ�ă����5�[�7y2`�e~�}�#� n���W�Y,(f��4�`BZ*n1�as�ϖ�����`�"��J������}��^ 1Њ}�_Ϟ:��aUŉ���e���ɗ�Ll���:Z�+�ꪭ�q�E���|�^�Qo%`����6ѓK�����:���27^`�y9Ƒ�ɛ�ן����XI��8e�u�kPc8/�S��,�	9# ��R�ihv?����MMS�+i8]cm�/��%���!F�'H�T�T.*Ȝ�*��QK��2��mM��Ϙ��W$���w�uBC�����LLQ�«jH�|����7u�*"&�Nu�)��_�<k�|ϯ